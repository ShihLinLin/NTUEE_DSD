module HA(A, B, S, C);
    input  A, B;
    output S, C;

    assign S = A ^ B;
    assign C = A & B;
endmodule

module FA(A, B, Cin, S, Cout);
    input  A, B, Cin;
    output S, Cout;

    assign S = A ^ B ^ Cin;
    assign Cout = (A & B) | (B & Cin) | (A & Cin);
    // assign Cout = (A & B) | (Cin & (A ^ B));
endmodule

module dadda (A, B, C);
    input  [31:0] A, B;
    output [31:0] C;
    
    // reg  [31:0] A, B, C_r;
    // wire [31:0] C;

    // assign C = C_r;

    wire s_1_1_8, s_1_2_8, s_1_3_8, s_1_4_8, s_1_5_8, s_1_6_8, s_1_7_8, s_1_8_8, s_1_9_8, s_1_10_8, s_1_11_8, s_1_12_8, s_1_13_8, s_1_14_8, s_1_15_8, s_1_16_8, s_1_17_8, s_1_18_8, s_1_19_8, s_1_20_8, s_1_21_8, s_1_22_8, s_1_23_8, s_1_24_8, s_1_25_8, s_1_26_8, s_1_27_8, s_1_28_8, s_1_29_8, s_1_30_8, s_1_31_8, s_1_32_8, s_2_2_8, s_2_3_8, s_2_4_8, s_2_5_8, s_2_6_8, s_2_7_8, s_2_8_8, s_2_9_8, s_2_10_8, s_2_11_8, s_2_12_8, s_2_13_8, s_2_14_8, s_2_15_8, s_2_16_8, s_2_17_8, s_2_18_8, s_2_19_8, s_2_20_8, s_2_21_8, s_2_22_8, s_2_23_8, s_2_24_8, s_2_25_8, s_2_26_8, s_2_27_8, s_2_28_8, s_2_29_8, s_2_30_8, s_2_31_8, s_2_32_8, s_3_3_8, s_3_4_8, s_3_5_8, s_3_6_8, s_3_7_8, s_3_8_8, s_3_9_8, s_3_10_8, s_3_11_8, s_3_12_8, s_3_13_8, s_3_14_8, s_3_15_8, s_3_16_8, s_3_17_8, s_3_18_8, s_3_19_8, s_3_20_8, s_3_21_8, s_3_22_8, s_3_23_8, s_3_24_8, s_3_25_8, s_3_26_8, s_3_27_8, s_3_28_8, s_3_29_8, s_3_30_8, s_3_31_8, s_3_32_8, s_4_4_8, s_4_5_8, s_4_6_8, s_4_7_8, s_4_8_8, s_4_9_8, s_4_10_8, s_4_11_8, s_4_12_8, s_4_13_8, s_4_14_8, s_4_15_8, s_4_16_8, s_4_17_8, s_4_18_8, s_4_19_8, s_4_20_8, s_4_21_8, s_4_22_8, s_4_23_8, s_4_24_8, s_4_25_8, s_4_26_8, s_4_27_8, s_4_28_8, s_4_29_8, s_4_30_8, s_4_31_8, s_4_32_8, s_5_5_8, s_5_6_8, s_5_7_8, s_5_8_8, s_5_9_8, s_5_10_8, s_5_11_8, s_5_12_8, s_5_13_8, s_5_14_8, s_5_15_8, s_5_16_8, s_5_17_8, s_5_18_8, s_5_19_8, s_5_20_8, s_5_21_8, s_5_22_8, s_5_23_8, s_5_24_8, s_5_25_8, s_5_26_8, s_5_27_8, s_5_28_8, s_5_29_8, s_5_30_8, s_5_31_8, s_5_32_8, s_6_6_8, s_6_7_8, s_6_8_8, s_6_9_8, s_6_10_8, s_6_11_8, s_6_12_8, s_6_13_8, s_6_14_8, s_6_15_8, s_6_16_8, s_6_17_8, s_6_18_8, s_6_19_8, s_6_20_8, s_6_21_8, s_6_22_8, s_6_23_8, s_6_24_8, s_6_25_8, s_6_26_8, s_6_27_8, s_6_28_8, s_6_29_8, s_6_30_8, s_6_31_8, s_6_32_8, s_7_7_8, s_7_8_8, s_7_9_8, s_7_10_8, s_7_11_8, s_7_12_8, s_7_13_8, s_7_14_8, s_7_15_8, s_7_16_8, s_7_17_8, s_7_18_8, s_7_19_8, s_7_20_8, s_7_21_8, s_7_22_8, s_7_23_8, s_7_24_8, s_7_25_8, s_7_26_8, s_7_27_8, s_7_28_8, s_7_29_8, s_7_30_8, s_7_31_8, s_7_32_8, s_8_8_8, s_8_9_8, s_8_10_8, s_8_11_8, s_8_12_8, s_8_13_8, s_8_14_8, s_8_15_8, s_8_16_8, s_8_17_8, s_8_18_8, s_8_19_8, s_8_20_8, s_8_21_8, s_8_22_8, s_8_23_8, s_8_24_8, s_8_25_8, s_8_26_8, s_8_27_8, s_8_28_8, s_8_29_8, s_8_30_8, s_8_31_8, s_8_32_8, s_9_9_8, s_9_10_8, s_9_11_8, s_9_12_8, s_9_13_8, s_9_14_8, s_9_15_8, s_9_16_8, s_9_17_8, s_9_18_8, s_9_19_8, s_9_20_8, s_9_21_8, s_9_22_8, s_9_23_8, s_9_24_8, s_9_25_8, s_9_26_8, s_9_27_8, s_9_28_8, s_9_29_8, s_9_30_8, s_9_31_8, s_9_32_8, s_10_10_8, s_10_11_8, s_10_12_8, s_10_13_8, s_10_14_8, s_10_15_8, s_10_16_8, s_10_17_8, s_10_18_8, s_10_19_8, s_10_20_8, s_10_21_8, s_10_22_8, s_10_23_8, s_10_24_8, s_10_25_8, s_10_26_8, s_10_27_8, s_10_28_8, s_10_29_8, s_10_30_8, s_10_31_8, s_10_32_8, s_11_11_8, s_11_12_8, s_11_13_8, s_11_14_8, s_11_15_8, s_11_16_8, s_11_17_8, s_11_18_8, s_11_19_8, s_11_20_8, s_11_21_8, s_11_22_8, s_11_23_8, s_11_24_8, s_11_25_8, s_11_26_8, s_11_27_8, s_11_28_8, s_11_29_8, s_11_30_8, s_11_31_8, s_11_32_8, s_12_12_8, s_12_13_8, s_12_14_8, s_12_15_8, s_12_16_8, s_12_17_8, s_12_18_8, s_12_19_8, s_12_20_8, s_12_21_8, s_12_22_8, s_12_23_8, s_12_24_8, s_12_25_8, s_12_26_8, s_12_27_8, s_12_28_8, s_12_29_8, s_12_30_8, s_12_31_8, s_12_32_8, s_13_13_8, s_13_14_8, s_13_15_8, s_13_16_8, s_13_17_8, s_13_18_8, s_13_19_8, s_13_20_8, s_13_21_8, s_13_22_8, s_13_23_8, s_13_24_8, s_13_25_8, s_13_26_8, s_13_27_8, s_13_28_8, s_13_29_8, s_13_30_8, s_13_31_8, s_13_32_8, s_14_14_8, s_14_15_8, s_14_16_8, s_14_17_8, s_14_18_8, s_14_19_8, s_14_20_8, s_14_21_8, s_14_22_8, s_14_23_8, s_14_24_8, s_14_25_8, s_14_26_8, s_14_27_8, s_14_28_8, s_14_29_8, s_14_30_8, s_14_31_8, s_14_32_8, s_15_15_8, s_15_16_8, s_15_17_8, s_15_18_8, s_15_19_8, s_15_20_8, s_15_21_8, s_15_22_8, s_15_23_8, s_15_24_8, s_15_25_8, s_15_26_8, s_15_27_8, s_15_28_8, s_15_29_8, s_15_30_8, s_15_31_8, s_15_32_8, s_16_16_8, s_16_17_8, s_16_18_8, s_16_19_8, s_16_20_8, s_16_21_8, s_16_22_8, s_16_23_8, s_16_24_8, s_16_25_8, s_16_26_8, s_16_27_8, s_16_28_8, s_16_29_8, s_16_30_8, s_16_31_8, s_16_32_8, s_17_17_8, s_17_18_8, s_17_19_8, s_17_20_8, s_17_21_8, s_17_22_8, s_17_23_8, s_17_24_8, s_17_25_8, s_17_26_8, s_17_27_8, s_17_28_8, s_17_29_8, s_17_30_8, s_17_31_8, s_17_32_8, s_18_18_8, s_18_19_8, s_18_20_8, s_18_21_8, s_18_22_8, s_18_23_8, s_18_24_8, s_18_25_8, s_18_26_8, s_18_27_8, s_18_28_8, s_18_29_8, s_18_30_8, s_18_31_8, s_18_32_8, s_19_19_8, s_19_20_8, s_19_21_8, s_19_22_8, s_19_23_8, s_19_24_8, s_19_25_8, s_19_26_8, s_19_27_8, s_19_28_8, s_19_29_8, s_19_30_8, s_19_31_8, s_19_32_8, s_20_20_8, s_20_21_8, s_20_22_8, s_20_23_8, s_20_24_8, s_20_25_8, s_20_26_8, s_20_27_8, s_20_28_8, s_20_29_8, s_20_30_8, s_20_31_8, s_20_32_8, s_21_21_8, s_21_22_8, s_21_23_8, s_21_24_8, s_21_25_8, s_21_26_8, s_21_27_8, s_21_28_8, s_21_29_8, s_21_30_8, s_21_31_8, s_21_32_8, s_22_22_8, s_22_23_8, s_22_24_8, s_22_25_8, s_22_26_8, s_22_27_8, s_22_28_8, s_22_29_8, s_22_30_8, s_22_31_8, s_22_32_8, s_23_23_8, s_23_24_8, s_23_25_8, s_23_26_8, s_23_27_8, s_23_28_8, s_23_29_8, s_23_30_8, s_23_31_8, s_23_32_8, s_24_24_8, s_24_25_8, s_24_26_8, s_24_27_8, s_24_28_8, s_24_29_8, s_24_30_8, s_24_31_8, s_24_32_8, s_25_25_8, s_25_26_8, s_25_27_8, s_25_28_8, s_25_29_8, s_25_30_8, s_25_31_8, s_25_32_8, s_26_26_8, s_26_27_8, s_26_28_8, s_26_29_8, s_26_30_8, s_26_31_8, s_26_32_8, s_27_27_8, s_27_28_8, s_27_29_8, s_27_30_8, s_27_31_8, s_27_32_8, s_28_28_8, s_28_29_8, s_28_30_8, s_28_31_8, s_28_32_8, s_29_29_8, s_29_30_8, s_29_31_8, s_29_32_8, s_30_30_8, s_30_31_8, s_30_32_8, s_31_31_8, s_31_32_8, s_32_32_8;
        wire s_1_1_7, s_2_2_7, s_1_2_7, s_3_3_7, s_2_3_7, s_1_3_7, s_4_4_7, s_3_4_7, s_2_4_7, s_1_4_7, s_5_5_7, s_4_5_7, s_3_5_7, s_2_5_7, s_1_5_7, s_6_6_7, s_5_6_7, s_4_6_7, s_3_6_7, s_2_6_7, s_1_6_7, s_7_7_7, s_6_7_7, s_5_7_7, s_4_7_7, s_3_7_7, s_2_7_7, s_1_7_7, s_8_8_7, s_7_8_7, s_6_8_7, s_5_8_7, s_4_8_7, s_3_8_7, s_2_8_7, s_1_8_7, s_9_9_7, s_8_9_7, s_7_9_7, s_6_9_7, s_5_9_7, s_4_9_7, s_3_9_7, s_2_9_7, s_1_9_7, s_10_10_7, s_9_10_7, s_8_10_7, s_7_10_7, s_6_10_7, s_5_10_7, s_4_10_7, s_3_10_7, s_2_10_7, s_1_10_7, s_11_11_7, s_10_11_7, s_9_11_7, s_8_11_7, s_7_11_7, s_6_11_7, s_5_11_7, s_4_11_7, s_3_11_7, s_2_11_7, s_1_11_7, s_12_12_7, s_11_12_7, s_10_12_7, s_9_12_7, s_8_12_7, s_7_12_7, s_6_12_7, s_5_12_7, s_4_12_7, s_3_12_7, s_2_12_7, s_1_12_7, s_13_13_7, s_12_13_7, s_11_13_7, s_10_13_7, s_9_13_7, s_8_13_7, s_7_13_7, s_6_13_7, s_5_13_7, s_4_13_7, s_3_13_7, s_2_13_7, s_1_13_7, s_14_14_7, s_13_14_7, s_12_14_7, s_11_14_7, s_10_14_7, s_9_14_7, s_8_14_7, s_7_14_7, s_6_14_7, s_5_14_7, s_4_14_7, s_3_14_7, s_2_14_7, s_1_14_7, s_15_15_7, s_14_15_7, s_13_15_7, s_12_15_7, s_11_15_7, s_10_15_7, s_9_15_7, s_8_15_7, s_7_15_7, s_6_15_7, s_5_15_7, s_4_15_7, s_3_15_7, s_2_15_7, s_1_15_7, s_16_16_7, s_15_16_7, s_14_16_7, s_13_16_7, s_12_16_7, s_11_16_7, s_10_16_7, s_9_16_7, s_8_16_7, s_7_16_7, s_6_16_7, s_5_16_7, s_4_16_7, s_3_16_7, s_2_16_7, s_1_16_7, s_17_17_7, s_16_17_7, s_15_17_7, s_14_17_7, s_13_17_7, s_12_17_7, s_11_17_7, s_10_17_7, s_9_17_7, s_8_17_7, s_7_17_7, s_6_17_7, s_5_17_7, s_4_17_7, s_3_17_7, s_2_17_7, s_1_17_7, s_18_18_7, s_17_18_7, s_16_18_7, s_15_18_7, s_14_18_7, s_13_18_7, s_12_18_7, s_11_18_7, s_10_18_7, s_9_18_7, s_8_18_7, s_7_18_7, s_6_18_7, s_5_18_7, s_4_18_7, s_3_18_7, s_2_18_7, s_1_18_7, s_19_19_7, s_18_19_7, s_17_19_7, s_16_19_7, s_15_19_7, s_14_19_7, s_13_19_7, s_12_19_7, s_11_19_7, s_10_19_7, s_9_19_7, s_8_19_7, s_7_19_7, s_6_19_7, s_5_19_7, s_4_19_7, s_3_19_7, s_2_19_7, s_1_19_7, s_20_20_7, s_19_20_7, s_18_20_7, s_17_20_7, s_16_20_7, s_15_20_7, s_14_20_7, s_13_20_7, s_12_20_7, s_11_20_7, s_10_20_7, s_9_20_7, s_8_20_7, s_7_20_7, s_6_20_7, s_5_20_7, s_4_20_7, s_3_20_7, s_2_20_7, s_1_20_7, s_21_21_7, s_20_21_7, s_19_21_7, s_18_21_7, s_17_21_7, s_16_21_7, s_15_21_7, s_14_21_7, s_13_21_7, s_12_21_7, s_11_21_7, s_10_21_7, s_9_21_7, s_8_21_7, s_7_21_7, s_6_21_7, s_5_21_7, s_4_21_7, s_3_21_7, s_2_21_7, s_1_21_7, s_22_22_7, s_21_22_7, s_20_22_7, s_19_22_7, s_18_22_7, s_17_22_7, s_16_22_7, s_15_22_7, s_14_22_7, s_13_22_7, s_12_22_7, s_11_22_7, s_10_22_7, s_9_22_7, s_8_22_7, s_7_22_7, s_6_22_7, s_5_22_7, s_4_22_7, s_3_22_7, s_2_22_7, s_1_22_7, s_23_23_7, s_22_23_7, s_21_23_7, s_20_23_7, s_19_23_7, s_18_23_7, s_17_23_7, s_16_23_7, s_15_23_7, s_14_23_7, s_13_23_7, s_12_23_7, s_11_23_7, s_10_23_7, s_9_23_7, s_8_23_7, s_7_23_7, s_6_23_7, s_5_23_7, s_4_23_7, s_3_23_7, s_2_23_7, s_1_23_7, s_24_24_7, s_23_24_7, s_22_24_7, s_21_24_7, s_20_24_7, s_19_24_7, s_18_24_7, s_17_24_7, s_16_24_7, s_15_24_7, s_14_24_7, s_13_24_7, s_12_24_7, s_11_24_7, s_10_24_7, s_9_24_7, s_8_24_7, s_7_24_7, s_6_24_7, s_5_24_7, s_4_24_7, s_3_24_7, s_2_24_7, s_1_24_7, s_25_25_7, s_24_25_7, s_23_25_7, s_22_25_7, s_21_25_7, s_20_25_7, s_19_25_7, s_18_25_7, s_17_25_7, s_16_25_7, s_15_25_7, s_14_25_7, s_13_25_7, s_12_25_7, s_11_25_7, s_10_25_7, s_9_25_7, s_8_25_7, s_7_25_7, s_6_25_7, s_5_25_7, s_4_25_7, s_3_25_7, s_2_25_7, s_1_25_7, s_26_26_7, s_25_26_7, s_24_26_7, s_23_26_7, s_22_26_7, s_21_26_7, s_20_26_7, s_19_26_7, s_18_26_7, s_17_26_7, s_16_26_7, s_15_26_7, s_14_26_7, s_13_26_7, s_12_26_7, s_11_26_7, s_10_26_7, s_9_26_7, s_8_26_7, s_7_26_7, s_6_26_7, s_5_26_7, s_4_26_7, s_3_26_7, s_2_26_7, s_1_26_7, s_27_27_7, s_26_27_7, s_25_27_7, s_24_27_7, s_23_27_7, s_22_27_7, s_21_27_7, s_20_27_7, s_19_27_7, s_18_27_7, s_17_27_7, s_16_27_7, s_15_27_7, s_14_27_7, s_13_27_7, s_12_27_7, s_11_27_7, s_10_27_7, s_9_27_7, s_8_27_7, s_7_27_7, s_6_27_7, s_5_27_7, s_4_27_7, s_3_27_7, s_2_27_7, s_1_27_7, s_28_28_7, s_27_28_7, s_26_28_7, s_25_28_7, s_24_28_7, s_23_28_7, s_22_28_7, s_21_28_7, s_20_28_7, s_19_28_7, s_18_28_7, s_17_28_7, s_16_28_7, s_15_28_7, s_14_28_7, s_13_28_7, s_12_28_7, s_11_28_7, s_10_28_7, s_9_28_7, s_8_28_7, s_7_28_7, s_6_28_7, s_5_28_7, s_4_28_7, s_3_28_7, s_2_28_7, s_1_28_7; 
    wire s_28_29_7, s_28_30_7; 
    wire s_27_29_7, s_26_29_7, s_25_29_7, s_24_29_7, s_23_29_7, s_22_29_7, s_21_29_7, s_20_29_7, s_19_29_7, s_18_29_7, s_17_29_7, s_16_29_7, s_15_29_7, s_14_29_7, s_13_29_7, s_12_29_7, s_11_29_7, s_10_29_7, s_9_29_7, s_8_29_7, s_7_29_7, s_6_29_7, s_5_29_7, s_4_29_7, s_3_29_7, s_2_29_7, s_1_29_7; 
    wire s_27_30_7, s_28_31_7; 
    wire s_26_30_7, s_27_31_7; 
    wire s_25_30_7, s_24_30_7, s_23_30_7, s_22_30_7, s_21_30_7, s_20_30_7, s_19_30_7, s_18_30_7, s_17_30_7, s_16_30_7, s_15_30_7, s_14_30_7, s_13_30_7, s_12_30_7, s_11_30_7, s_10_30_7, s_9_30_7, s_8_30_7, s_7_30_7, s_6_30_7, s_5_30_7, s_4_30_7, s_3_30_7, s_2_30_7, s_1_30_7; 
    wire s_26_31_7, s_28_32_7; 
    wire s_25_31_7, s_27_32_7; 
    wire s_24_31_7, s_26_32_7; 
    wire s_23_31_7, s_22_31_7, s_21_31_7, s_20_31_7, s_19_31_7, s_18_31_7, s_17_31_7, s_16_31_7, s_15_31_7, s_14_31_7, s_13_31_7, s_12_31_7, s_11_31_7, s_10_31_7, s_9_31_7, s_8_31_7, s_7_31_7, s_6_31_7, s_5_31_7, s_4_31_7, s_3_31_7, s_2_31_7, s_1_31_7; 
    wire s_25_32_7, s_28_33_7; 
    wire s_24_32_7, s_27_33_7; 
    wire s_23_32_7, s_26_33_7; 
    wire s_22_32_7, s_25_33_7; 
    wire s_21_32_7, s_20_32_7, s_19_32_7, s_18_32_7, s_17_32_7, s_16_32_7, s_15_32_7, s_14_32_7, s_13_32_7, s_12_32_7, s_11_32_7, s_10_32_7, s_9_32_7, s_8_32_7, s_7_32_7, s_6_32_7, s_5_32_7, s_4_32_7, s_3_32_7, s_2_32_7, s_1_32_7; 
    // total 4 half adders and 6 full adders
    // d_8 = 28 done

    wire s_1_1_6, s_2_2_6, s_1_2_6, s_3_3_6, s_2_3_6, s_1_3_6, s_4_4_6, s_3_4_6, s_2_4_6, s_1_4_6, s_5_5_6, s_4_5_6, s_3_5_6, s_2_5_6, s_1_5_6, s_6_6_6, s_5_6_6, s_4_6_6, s_3_6_6, s_2_6_6, s_1_6_6, s_7_7_6, s_6_7_6, s_5_7_6, s_4_7_6, s_3_7_6, s_2_7_6, s_1_7_6, s_8_8_6, s_7_8_6, s_6_8_6, s_5_8_6, s_4_8_6, s_3_8_6, s_2_8_6, s_1_8_6, s_9_9_6, s_8_9_6, s_7_9_6, s_6_9_6, s_5_9_6, s_4_9_6, s_3_9_6, s_2_9_6, s_1_9_6, s_10_10_6, s_9_10_6, s_8_10_6, s_7_10_6, s_6_10_6, s_5_10_6, s_4_10_6, s_3_10_6, s_2_10_6, s_1_10_6, s_11_11_6, s_10_11_6, s_9_11_6, s_8_11_6, s_7_11_6, s_6_11_6, s_5_11_6, s_4_11_6, s_3_11_6, s_2_11_6, s_1_11_6, s_12_12_6, s_11_12_6, s_10_12_6, s_9_12_6, s_8_12_6, s_7_12_6, s_6_12_6, s_5_12_6, s_4_12_6, s_3_12_6, s_2_12_6, s_1_12_6, s_13_13_6, s_12_13_6, s_11_13_6, s_10_13_6, s_9_13_6, s_8_13_6, s_7_13_6, s_6_13_6, s_5_13_6, s_4_13_6, s_3_13_6, s_2_13_6, s_1_13_6, s_14_14_6, s_13_14_6, s_12_14_6, s_11_14_6, s_10_14_6, s_9_14_6, s_8_14_6, s_7_14_6, s_6_14_6, s_5_14_6, s_4_14_6, s_3_14_6, s_2_14_6, s_1_14_6, s_15_15_6, s_14_15_6, s_13_15_6, s_12_15_6, s_11_15_6, s_10_15_6, s_9_15_6, s_8_15_6, s_7_15_6, s_6_15_6, s_5_15_6, s_4_15_6, s_3_15_6, s_2_15_6, s_1_15_6, s_16_16_6, s_15_16_6, s_14_16_6, s_13_16_6, s_12_16_6, s_11_16_6, s_10_16_6, s_9_16_6, s_8_16_6, s_7_16_6, s_6_16_6, s_5_16_6, s_4_16_6, s_3_16_6, s_2_16_6, s_1_16_6, s_17_17_6, s_16_17_6, s_15_17_6, s_14_17_6, s_13_17_6, s_12_17_6, s_11_17_6, s_10_17_6, s_9_17_6, s_8_17_6, s_7_17_6, s_6_17_6, s_5_17_6, s_4_17_6, s_3_17_6, s_2_17_6, s_1_17_6, s_18_18_6, s_17_18_6, s_16_18_6, s_15_18_6, s_14_18_6, s_13_18_6, s_12_18_6, s_11_18_6, s_10_18_6, s_9_18_6, s_8_18_6, s_7_18_6, s_6_18_6, s_5_18_6, s_4_18_6, s_3_18_6, s_2_18_6, s_1_18_6, s_19_19_6, s_18_19_6, s_17_19_6, s_16_19_6, s_15_19_6, s_14_19_6, s_13_19_6, s_12_19_6, s_11_19_6, s_10_19_6, s_9_19_6, s_8_19_6, s_7_19_6, s_6_19_6, s_5_19_6, s_4_19_6, s_3_19_6, s_2_19_6, s_1_19_6; 
    wire s_19_20_6, s_19_21_6; 
    wire s_18_20_6, s_17_20_6, s_16_20_6, s_15_20_6, s_14_20_6, s_13_20_6, s_12_20_6, s_11_20_6, s_10_20_6, s_9_20_6, s_8_20_6, s_7_20_6, s_6_20_6, s_5_20_6, s_4_20_6, s_3_20_6, s_2_20_6, s_1_20_6; 
    wire s_18_21_6, s_19_22_6; 
    wire s_17_21_6, s_18_22_6; 
    wire s_16_21_6, s_15_21_6, s_14_21_6, s_13_21_6, s_12_21_6, s_11_21_6, s_10_21_6, s_9_21_6, s_8_21_6, s_7_21_6, s_6_21_6, s_5_21_6, s_4_21_6, s_3_21_6, s_2_21_6, s_1_21_6; 
    wire s_17_22_6, s_19_23_6; 
    wire s_16_22_6, s_18_23_6; 
    wire s_15_22_6, s_17_23_6; 
    wire s_14_22_6, s_13_22_6, s_12_22_6, s_11_22_6, s_10_22_6, s_9_22_6, s_8_22_6, s_7_22_6, s_6_22_6, s_5_22_6, s_4_22_6, s_3_22_6, s_2_22_6, s_1_22_6; 
    wire s_16_23_6, s_19_24_6; 
    wire s_15_23_6, s_18_24_6; 
    wire s_14_23_6, s_17_24_6; 
    wire s_13_23_6, s_16_24_6; 
    wire s_12_23_6, s_11_23_6, s_10_23_6, s_9_23_6, s_8_23_6, s_7_23_6, s_6_23_6, s_5_23_6, s_4_23_6, s_3_23_6, s_2_23_6, s_1_23_6; 
    wire s_15_24_6, s_19_25_6; 
    wire s_14_24_6, s_18_25_6; 
    wire s_13_24_6, s_17_25_6; 
    wire s_12_24_6, s_16_25_6; 
    wire s_11_24_6, s_15_25_6; 
    wire s_10_24_6, s_9_24_6, s_8_24_6, s_7_24_6, s_6_24_6, s_5_24_6, s_4_24_6, s_3_24_6, s_2_24_6, s_1_24_6; 
    wire s_14_25_6, s_19_26_6; 
    wire s_13_25_6, s_18_26_6; 
    wire s_12_25_6, s_17_26_6; 
    wire s_11_25_6, s_16_26_6; 
    wire s_10_25_6, s_15_26_6; 
    wire s_9_25_6, s_14_26_6; 
    wire s_8_25_6, s_7_25_6, s_6_25_6, s_5_25_6, s_4_25_6, s_3_25_6, s_2_25_6, s_1_25_6; 
    wire s_13_26_6, s_19_27_6; 
    wire s_12_26_6, s_18_27_6; 
    wire s_11_26_6, s_17_27_6; 
    wire s_10_26_6, s_16_27_6; 
    wire s_9_26_6, s_15_27_6; 
    wire s_8_26_6, s_14_27_6; 
    wire s_7_26_6, s_13_27_6; 
    wire s_6_26_6, s_5_26_6, s_4_26_6, s_3_26_6, s_2_26_6, s_1_26_6; 
    wire s_12_27_6, s_19_28_6; 
    wire s_11_27_6, s_18_28_6; 
    wire s_10_27_6, s_17_28_6; 
    wire s_9_27_6, s_16_28_6; 
    wire s_8_27_6, s_15_28_6; 
    wire s_7_27_6, s_14_28_6; 
    wire s_6_27_6, s_13_28_6; 
    wire s_5_27_6, s_12_28_6; 
    wire s_4_27_6, s_3_27_6, s_2_27_6, s_1_27_6; 
    wire s_11_28_6, s_19_29_6; 
    wire s_10_28_6, s_18_29_6; 
    wire s_9_28_6, s_17_29_6; 
    wire s_8_28_6, s_16_29_6; 
    wire s_7_28_6, s_15_29_6; 
    wire s_6_28_6, s_14_29_6; 
    wire s_5_28_6, s_13_29_6; 
    wire s_4_28_6, s_12_29_6; 
    wire s_3_28_6, s_11_29_6; 
    wire s_2_28_6, s_1_28_6; 
    wire s_10_29_6, s_19_30_6; 
    wire s_9_29_6, s_18_30_6; 
    wire s_8_29_6, s_17_30_6; 
    wire s_7_29_6, s_16_30_6; 
    wire s_6_29_6, s_15_30_6; 
    wire s_5_29_6, s_14_30_6; 
    wire s_4_29_6, s_13_30_6; 
    wire s_3_29_6, s_12_30_6; 
    wire s_2_29_6, s_11_30_6; 
    wire s_1_29_6; 
    wire s_10_30_6, s_19_31_6; 
    wire s_9_30_6, s_18_31_6; 
    wire s_8_30_6, s_17_31_6; 
    wire s_7_30_6, s_16_31_6; 
    wire s_6_30_6, s_15_31_6; 
    wire s_5_30_6, s_14_31_6; 
    wire s_4_30_6, s_13_31_6; 
    wire s_3_30_6, s_12_31_6; 
    wire s_2_30_6, s_11_31_6; 
    wire s_1_30_6; 
    wire s_10_31_6, s_19_32_6; 
    wire s_9_31_6, s_18_32_6; 
    wire s_8_31_6, s_17_32_6; 
    wire s_7_31_6, s_16_32_6; 
    wire s_6_31_6, s_15_32_6; 
    wire s_5_31_6, s_14_32_6; 
    wire s_4_31_6, s_13_32_6; 
    wire s_3_31_6, s_12_32_6; 
    wire s_2_31_6, s_11_32_6; 
    wire s_1_31_6; 
    wire s_10_32_6, s_19_33_6; 
    wire s_9_32_6, s_18_33_6; 
    wire s_8_32_6, s_17_33_6; 
    wire s_7_32_6, s_16_33_6; 
    wire s_6_32_6, s_15_33_6; 
    wire s_5_32_6, s_14_33_6; 
    wire s_4_32_6, s_13_33_6; 
    wire s_3_32_6, s_12_33_6; 
    wire s_2_32_6, s_11_33_6; 
    wire s_1_32_6; 
    // total 9 half adders and 72 full adders
    // d_7 = 19 done

    wire s_1_1_5, s_2_2_5, s_1_2_5, s_3_3_5, s_2_3_5, s_1_3_5, s_4_4_5, s_3_4_5, s_2_4_5, s_1_4_5, s_5_5_5, s_4_5_5, s_3_5_5, s_2_5_5, s_1_5_5, s_6_6_5, s_5_6_5, s_4_6_5, s_3_6_5, s_2_6_5, s_1_6_5, s_7_7_5, s_6_7_5, s_5_7_5, s_4_7_5, s_3_7_5, s_2_7_5, s_1_7_5, s_8_8_5, s_7_8_5, s_6_8_5, s_5_8_5, s_4_8_5, s_3_8_5, s_2_8_5, s_1_8_5, s_9_9_5, s_8_9_5, s_7_9_5, s_6_9_5, s_5_9_5, s_4_9_5, s_3_9_5, s_2_9_5, s_1_9_5, s_10_10_5, s_9_10_5, s_8_10_5, s_7_10_5, s_6_10_5, s_5_10_5, s_4_10_5, s_3_10_5, s_2_10_5, s_1_10_5, s_11_11_5, s_10_11_5, s_9_11_5, s_8_11_5, s_7_11_5, s_6_11_5, s_5_11_5, s_4_11_5, s_3_11_5, s_2_11_5, s_1_11_5, s_12_12_5, s_11_12_5, s_10_12_5, s_9_12_5, s_8_12_5, s_7_12_5, s_6_12_5, s_5_12_5, s_4_12_5, s_3_12_5, s_2_12_5, s_1_12_5, s_13_13_5, s_12_13_5, s_11_13_5, s_10_13_5, s_9_13_5, s_8_13_5, s_7_13_5, s_6_13_5, s_5_13_5, s_4_13_5, s_3_13_5, s_2_13_5, s_1_13_5; 
    wire s_13_14_5, s_13_15_5; 
    wire s_12_14_5, s_11_14_5, s_10_14_5, s_9_14_5, s_8_14_5, s_7_14_5, s_6_14_5, s_5_14_5, s_4_14_5, s_3_14_5, s_2_14_5, s_1_14_5; 
    wire s_12_15_5, s_13_16_5; 
    wire s_11_15_5, s_12_16_5; 
    wire s_10_15_5, s_9_15_5, s_8_15_5, s_7_15_5, s_6_15_5, s_5_15_5, s_4_15_5, s_3_15_5, s_2_15_5, s_1_15_5; 
    wire s_11_16_5, s_13_17_5; 
    wire s_10_16_5, s_12_17_5; 
    wire s_9_16_5, s_11_17_5; 
    wire s_8_16_5, s_7_16_5, s_6_16_5, s_5_16_5, s_4_16_5, s_3_16_5, s_2_16_5, s_1_16_5; 
    wire s_10_17_5, s_13_18_5; 
    wire s_9_17_5, s_12_18_5; 
    wire s_8_17_5, s_11_18_5; 
    wire s_7_17_5, s_10_18_5; 
    wire s_6_17_5, s_5_17_5, s_4_17_5, s_3_17_5, s_2_17_5, s_1_17_5; 
    wire s_9_18_5, s_13_19_5; 
    wire s_8_18_5, s_12_19_5; 
    wire s_7_18_5, s_11_19_5; 
    wire s_6_18_5, s_10_19_5; 
    wire s_5_18_5, s_9_19_5; 
    wire s_4_18_5, s_3_18_5, s_2_18_5, s_1_18_5; 
    wire s_8_19_5, s_13_20_5; 
    wire s_7_19_5, s_12_20_5; 
    wire s_6_19_5, s_11_20_5; 
    wire s_5_19_5, s_10_20_5; 
    wire s_4_19_5, s_9_20_5; 
    wire s_3_19_5, s_8_20_5; 
    wire s_2_19_5, s_1_19_5; 
    wire s_7_20_5, s_13_21_5; 
    wire s_6_20_5, s_12_21_5; 
    wire s_5_20_5, s_11_21_5; 
    wire s_4_20_5, s_10_21_5; 
    wire s_3_20_5, s_9_21_5; 
    wire s_2_20_5, s_8_21_5; 
    wire s_1_20_5; 
    wire s_7_21_5, s_13_22_5; 
    wire s_6_21_5, s_12_22_5; 
    wire s_5_21_5, s_11_22_5; 
    wire s_4_21_5, s_10_22_5; 
    wire s_3_21_5, s_9_22_5; 
    wire s_2_21_5, s_8_22_5; 
    wire s_1_21_5; 
    wire s_7_22_5, s_13_23_5; 
    wire s_6_22_5, s_12_23_5; 
    wire s_5_22_5, s_11_23_5; 
    wire s_4_22_5, s_10_23_5; 
    wire s_3_22_5, s_9_23_5; 
    wire s_2_22_5, s_8_23_5; 
    wire s_1_22_5; 
    wire s_7_23_5, s_13_24_5; 
    wire s_6_23_5, s_12_24_5; 
    wire s_5_23_5, s_11_24_5; 
    wire s_4_23_5, s_10_24_5; 
    wire s_3_23_5, s_9_24_5; 
    wire s_2_23_5, s_8_24_5; 
    wire s_1_23_5; 
    wire s_7_24_5, s_13_25_5; 
    wire s_6_24_5, s_12_25_5; 
    wire s_5_24_5, s_11_25_5; 
    wire s_4_24_5, s_10_25_5; 
    wire s_3_24_5, s_9_25_5; 
    wire s_2_24_5, s_8_25_5; 
    wire s_1_24_5; 
    wire s_7_25_5, s_13_26_5; 
    wire s_6_25_5, s_12_26_5; 
    wire s_5_25_5, s_11_26_5; 
    wire s_4_25_5, s_10_26_5; 
    wire s_3_25_5, s_9_26_5; 
    wire s_2_25_5, s_8_26_5; 
    wire s_1_25_5; 
    wire s_7_26_5, s_13_27_5; 
    wire s_6_26_5, s_12_27_5; 
    wire s_5_26_5, s_11_27_5; 
    wire s_4_26_5, s_10_27_5; 
    wire s_3_26_5, s_9_27_5; 
    wire s_2_26_5, s_8_27_5; 
    wire s_1_26_5; 
    wire s_7_27_5, s_13_28_5; 
    wire s_6_27_5, s_12_28_5; 
    wire s_5_27_5, s_11_28_5; 
    wire s_4_27_5, s_10_28_5; 
    wire s_3_27_5, s_9_28_5; 
    wire s_2_27_5, s_8_28_5; 
    wire s_1_27_5; 
    wire s_7_28_5, s_13_29_5; 
    wire s_6_28_5, s_12_29_5; 
    wire s_5_28_5, s_11_29_5; 
    wire s_4_28_5, s_10_29_5; 
    wire s_3_28_5, s_9_29_5; 
    wire s_2_28_5, s_8_29_5; 
    wire s_1_28_5; 
    wire s_7_29_5, s_13_30_5; 
    wire s_6_29_5, s_12_30_5; 
    wire s_5_29_5, s_11_30_5; 
    wire s_4_29_5, s_10_30_5; 
    wire s_3_29_5, s_9_30_5; 
    wire s_2_29_5, s_8_30_5; 
    wire s_1_29_5; 
    wire s_7_30_5, s_13_31_5; 
    wire s_6_30_5, s_12_31_5; 
    wire s_5_30_5, s_11_31_5; 
    wire s_4_30_5, s_10_31_5; 
    wire s_3_30_5, s_9_31_5; 
    wire s_2_30_5, s_8_31_5; 
    wire s_1_30_5; 
    wire s_7_31_5, s_13_32_5; 
    wire s_6_31_5, s_12_32_5; 
    wire s_5_31_5, s_11_32_5; 
    wire s_4_31_5, s_10_32_5; 
    wire s_3_31_5, s_9_32_5; 
    wire s_2_31_5, s_8_32_5; 
    wire s_1_31_5; 
    wire s_7_32_5, s_13_33_5; 
    wire s_6_32_5, s_12_33_5; 
    wire s_5_32_5, s_11_33_5; 
    wire s_4_32_5, s_10_33_5; 
    wire s_3_32_5, s_9_33_5; 
    wire s_2_32_5, s_8_33_5; 
    wire s_1_32_5; 
    // total 6 half adders and 93 full adders
    // d_6 = 13 done

    wire s_1_1_4, s_2_2_4, s_1_2_4, s_3_3_4, s_2_3_4, s_1_3_4, s_4_4_4, s_3_4_4, s_2_4_4, s_1_4_4, s_5_5_4, s_4_5_4, s_3_5_4, s_2_5_4, s_1_5_4, s_6_6_4, s_5_6_4, s_4_6_4, s_3_6_4, s_2_6_4, s_1_6_4, s_7_7_4, s_6_7_4, s_5_7_4, s_4_7_4, s_3_7_4, s_2_7_4, s_1_7_4, s_8_8_4, s_7_8_4, s_6_8_4, s_5_8_4, s_4_8_4, s_3_8_4, s_2_8_4, s_1_8_4, s_9_9_4, s_8_9_4, s_7_9_4, s_6_9_4, s_5_9_4, s_4_9_4, s_3_9_4, s_2_9_4, s_1_9_4; 
    wire s_9_10_4, s_9_11_4; 
    wire s_8_10_4, s_7_10_4, s_6_10_4, s_5_10_4, s_4_10_4, s_3_10_4, s_2_10_4, s_1_10_4; 
    wire s_8_11_4, s_9_12_4; 
    wire s_7_11_4, s_8_12_4; 
    wire s_6_11_4, s_5_11_4, s_4_11_4, s_3_11_4, s_2_11_4, s_1_11_4; 
    wire s_7_12_4, s_9_13_4; 
    wire s_6_12_4, s_8_13_4; 
    wire s_5_12_4, s_7_13_4; 
    wire s_4_12_4, s_3_12_4, s_2_12_4, s_1_12_4; 
    wire s_6_13_4, s_9_14_4; 
    wire s_5_13_4, s_8_14_4; 
    wire s_4_13_4, s_7_14_4; 
    wire s_3_13_4, s_6_14_4; 
    wire s_2_13_4, s_1_13_4; 
    wire s_5_14_4, s_9_15_4; 
    wire s_4_14_4, s_8_15_4; 
    wire s_3_14_4, s_7_15_4; 
    wire s_2_14_4, s_6_15_4; 
    wire s_1_14_4; 
    wire s_5_15_4, s_9_16_4; 
    wire s_4_15_4, s_8_16_4; 
    wire s_3_15_4, s_7_16_4; 
    wire s_2_15_4, s_6_16_4; 
    wire s_1_15_4; 
    wire s_5_16_4, s_9_17_4; 
    wire s_4_16_4, s_8_17_4; 
    wire s_3_16_4, s_7_17_4; 
    wire s_2_16_4, s_6_17_4; 
    wire s_1_16_4; 
    wire s_5_17_4, s_9_18_4; 
    wire s_4_17_4, s_8_18_4; 
    wire s_3_17_4, s_7_18_4; 
    wire s_2_17_4, s_6_18_4; 
    wire s_1_17_4; 
    wire s_5_18_4, s_9_19_4; 
    wire s_4_18_4, s_8_19_4; 
    wire s_3_18_4, s_7_19_4; 
    wire s_2_18_4, s_6_19_4; 
    wire s_1_18_4; 
    wire s_5_19_4, s_9_20_4; 
    wire s_4_19_4, s_8_20_4; 
    wire s_3_19_4, s_7_20_4; 
    wire s_2_19_4, s_6_20_4; 
    wire s_1_19_4; 
    wire s_5_20_4, s_9_21_4; 
    wire s_4_20_4, s_8_21_4; 
    wire s_3_20_4, s_7_21_4; 
    wire s_2_20_4, s_6_21_4; 
    wire s_1_20_4; 
    wire s_5_21_4, s_9_22_4; 
    wire s_4_21_4, s_8_22_4; 
    wire s_3_21_4, s_7_22_4; 
    wire s_2_21_4, s_6_22_4; 
    wire s_1_21_4; 
    wire s_5_22_4, s_9_23_4; 
    wire s_4_22_4, s_8_23_4; 
    wire s_3_22_4, s_7_23_4; 
    wire s_2_22_4, s_6_23_4; 
    wire s_1_22_4; 
    wire s_5_23_4, s_9_24_4; 
    wire s_4_23_4, s_8_24_4; 
    wire s_3_23_4, s_7_24_4; 
    wire s_2_23_4, s_6_24_4; 
    wire s_1_23_4; 
    wire s_5_24_4, s_9_25_4; 
    wire s_4_24_4, s_8_25_4; 
    wire s_3_24_4, s_7_25_4; 
    wire s_2_24_4, s_6_25_4; 
    wire s_1_24_4; 
    wire s_5_25_4, s_9_26_4; 
    wire s_4_25_4, s_8_26_4; 
    wire s_3_25_4, s_7_26_4; 
    wire s_2_25_4, s_6_26_4; 
    wire s_1_25_4; 
    wire s_5_26_4, s_9_27_4; 
    wire s_4_26_4, s_8_27_4; 
    wire s_3_26_4, s_7_27_4; 
    wire s_2_26_4, s_6_27_4; 
    wire s_1_26_4; 
    wire s_5_27_4, s_9_28_4; 
    wire s_4_27_4, s_8_28_4; 
    wire s_3_27_4, s_7_28_4; 
    wire s_2_27_4, s_6_28_4; 
    wire s_1_27_4; 
    wire s_5_28_4, s_9_29_4; 
    wire s_4_28_4, s_8_29_4; 
    wire s_3_28_4, s_7_29_4; 
    wire s_2_28_4, s_6_29_4; 
    wire s_1_28_4; 
    wire s_5_29_4, s_9_30_4; 
    wire s_4_29_4, s_8_30_4; 
    wire s_3_29_4, s_7_30_4; 
    wire s_2_29_4, s_6_30_4; 
    wire s_1_29_4; 
    wire s_5_30_4, s_9_31_4; 
    wire s_4_30_4, s_8_31_4; 
    wire s_3_30_4, s_7_31_4; 
    wire s_2_30_4, s_6_31_4; 
    wire s_1_30_4; 
    wire s_5_31_4, s_9_32_4; 
    wire s_4_31_4, s_8_32_4; 
    wire s_3_31_4, s_7_32_4; 
    wire s_2_31_4, s_6_32_4; 
    wire s_1_31_4; 
    wire s_5_32_4, s_9_33_4; 
    wire s_4_32_4, s_8_33_4; 
    wire s_3_32_4, s_7_33_4; 
    wire s_2_32_4, s_6_33_4; 
    wire s_1_32_4; 
    // total 4 half adders and 82 full adders
    // d_5 = 9 done

    wire s_1_1_3, s_2_2_3, s_1_2_3, s_3_3_3, s_2_3_3, s_1_3_3, s_4_4_3, s_3_4_3, s_2_4_3, s_1_4_3, s_5_5_3, s_4_5_3, s_3_5_3, s_2_5_3, s_1_5_3, s_6_6_3, s_5_6_3, s_4_6_3, s_3_6_3, s_2_6_3, s_1_6_3; 
    wire s_6_7_3, s_6_8_3; 
    wire s_5_7_3, s_4_7_3, s_3_7_3, s_2_7_3, s_1_7_3; 
    wire s_5_8_3, s_6_9_3; 
    wire s_4_8_3, s_5_9_3; 
    wire s_3_8_3, s_2_8_3, s_1_8_3; 
    wire s_4_9_3, s_6_10_3; 
    wire s_3_9_3, s_5_10_3; 
    wire s_2_9_3, s_4_10_3; 
    wire s_1_9_3; 
    wire s_3_10_3, s_6_11_3; 
    wire s_2_10_3, s_5_11_3; 
    wire s_1_10_3, s_4_11_3; 
    wire s_3_11_3, s_6_12_3; 
    wire s_2_11_3, s_5_12_3; 
    wire s_1_11_3, s_4_12_3; 
    wire s_3_12_3, s_6_13_3; 
    wire s_2_12_3, s_5_13_3; 
    wire s_1_12_3, s_4_13_3; 
    wire s_3_13_3, s_6_14_3; 
    wire s_2_13_3, s_5_14_3; 
    wire s_1_13_3, s_4_14_3; 
    wire s_3_14_3, s_6_15_3; 
    wire s_2_14_3, s_5_15_3; 
    wire s_1_14_3, s_4_15_3; 
    wire s_3_15_3, s_6_16_3; 
    wire s_2_15_3, s_5_16_3; 
    wire s_1_15_3, s_4_16_3; 
    wire s_3_16_3, s_6_17_3; 
    wire s_2_16_3, s_5_17_3; 
    wire s_1_16_3, s_4_17_3; 
    wire s_3_17_3, s_6_18_3; 
    wire s_2_17_3, s_5_18_3; 
    wire s_1_17_3, s_4_18_3; 
    wire s_3_18_3, s_6_19_3; 
    wire s_2_18_3, s_5_19_3; 
    wire s_1_18_3, s_4_19_3; 
    wire s_3_19_3, s_6_20_3; 
    wire s_2_19_3, s_5_20_3; 
    wire s_1_19_3, s_4_20_3; 
    wire s_3_20_3, s_6_21_3; 
    wire s_2_20_3, s_5_21_3; 
    wire s_1_20_3, s_4_21_3; 
    wire s_3_21_3, s_6_22_3; 
    wire s_2_21_3, s_5_22_3; 
    wire s_1_21_3, s_4_22_3; 
    wire s_3_22_3, s_6_23_3; 
    wire s_2_22_3, s_5_23_3; 
    wire s_1_22_3, s_4_23_3; 
    wire s_3_23_3, s_6_24_3; 
    wire s_2_23_3, s_5_24_3; 
    wire s_1_23_3, s_4_24_3; 
    wire s_3_24_3, s_6_25_3; 
    wire s_2_24_3, s_5_25_3; 
    wire s_1_24_3, s_4_25_3; 
    wire s_3_25_3, s_6_26_3; 
    wire s_2_25_3, s_5_26_3; 
    wire s_1_25_3, s_4_26_3; 
    wire s_3_26_3, s_6_27_3; 
    wire s_2_26_3, s_5_27_3; 
    wire s_1_26_3, s_4_27_3; 
    wire s_3_27_3, s_6_28_3; 
    wire s_2_27_3, s_5_28_3; 
    wire s_1_27_3, s_4_28_3; 
    wire s_3_28_3, s_6_29_3; 
    wire s_2_28_3, s_5_29_3; 
    wire s_1_28_3, s_4_29_3; 
    wire s_3_29_3, s_6_30_3; 
    wire s_2_29_3, s_5_30_3; 
    wire s_1_29_3, s_4_30_3; 
    wire s_3_30_3, s_6_31_3; 
    wire s_2_30_3, s_5_31_3; 
    wire s_1_30_3, s_4_31_3; 
    wire s_3_31_3, s_6_32_3; 
    wire s_2_31_3, s_5_32_3; 
    wire s_1_31_3, s_4_32_3; 
    wire s_3_32_3, s_6_33_3; 
    wire s_2_32_3, s_5_33_3; 
    wire s_1_32_3, s_4_33_3; 
    // total 3 half adders and 72 full adders
    // d_4 = 6 done

    wire s_1_1_2, s_2_2_2, s_1_2_2, s_3_3_2, s_2_3_2, s_1_3_2, s_4_4_2, s_3_4_2, s_2_4_2, s_1_4_2; 
    wire s_4_5_2, s_4_6_2; 
    wire s_3_5_2, s_2_5_2, s_1_5_2; 
    wire s_3_6_2, s_4_7_2; 
    wire s_2_6_2, s_3_7_2; 
    wire s_1_6_2; 
    wire s_2_7_2, s_4_8_2; 
    wire s_1_7_2, s_3_8_2; 
    wire s_2_8_2, s_4_9_2; 
    wire s_1_8_2, s_3_9_2; 
    wire s_2_9_2, s_4_10_2; 
    wire s_1_9_2, s_3_10_2; 
    wire s_2_10_2, s_4_11_2; 
    wire s_1_10_2, s_3_11_2; 
    wire s_2_11_2, s_4_12_2; 
    wire s_1_11_2, s_3_12_2; 
    wire s_2_12_2, s_4_13_2; 
    wire s_1_12_2, s_3_13_2; 
    wire s_2_13_2, s_4_14_2; 
    wire s_1_13_2, s_3_14_2; 
    wire s_2_14_2, s_4_15_2; 
    wire s_1_14_2, s_3_15_2; 
    wire s_2_15_2, s_4_16_2; 
    wire s_1_15_2, s_3_16_2; 
    wire s_2_16_2, s_4_17_2; 
    wire s_1_16_2, s_3_17_2; 
    wire s_2_17_2, s_4_18_2; 
    wire s_1_17_2, s_3_18_2; 
    wire s_2_18_2, s_4_19_2; 
    wire s_1_18_2, s_3_19_2; 
    wire s_2_19_2, s_4_20_2; 
    wire s_1_19_2, s_3_20_2; 
    wire s_2_20_2, s_4_21_2; 
    wire s_1_20_2, s_3_21_2; 
    wire s_2_21_2, s_4_22_2; 
    wire s_1_21_2, s_3_22_2; 
    wire s_2_22_2, s_4_23_2; 
    wire s_1_22_2, s_3_23_2; 
    wire s_2_23_2, s_4_24_2; 
    wire s_1_23_2, s_3_24_2; 
    wire s_2_24_2, s_4_25_2; 
    wire s_1_24_2, s_3_25_2; 
    wire s_2_25_2, s_4_26_2; 
    wire s_1_25_2, s_3_26_2; 
    wire s_2_26_2, s_4_27_2; 
    wire s_1_26_2, s_3_27_2; 
    wire s_2_27_2, s_4_28_2; 
    wire s_1_27_2, s_3_28_2; 
    wire s_2_28_2, s_4_29_2; 
    wire s_1_28_2, s_3_29_2; 
    wire s_2_29_2, s_4_30_2; 
    wire s_1_29_2, s_3_30_2; 
    wire s_2_30_2, s_4_31_2; 
    wire s_1_30_2, s_3_31_2; 
    wire s_2_31_2, s_4_32_2; 
    wire s_1_31_2, s_3_32_2; 
    wire s_2_32_2, s_4_33_2; 
    wire s_1_32_2, s_3_33_2; 
    // total 2 half adders and 53 full adders
    // d_3 = 4 done

    wire s_1_1_1, s_2_2_1, s_1_2_1, s_3_3_1, s_2_3_1, s_1_3_1; 
    wire s_3_4_1, s_3_5_1; 
    wire s_2_4_1, s_1_4_1; 
    wire s_2_5_1, s_3_6_1; 
    wire s_1_5_1; 
    wire s_2_6_1, s_3_7_1; 
    wire s_1_6_1; 
    wire s_2_7_1, s_3_8_1; 
    wire s_1_7_1; 
    wire s_2_8_1, s_3_9_1; 
    wire s_1_8_1; 
    wire s_2_9_1, s_3_10_1; 
    wire s_1_9_1; 
    wire s_2_10_1, s_3_11_1; 
    wire s_1_10_1; 
    wire s_2_11_1, s_3_12_1; 
    wire s_1_11_1; 
    wire s_2_12_1, s_3_13_1; 
    wire s_1_12_1; 
    wire s_2_13_1, s_3_14_1; 
    wire s_1_13_1; 
    wire s_2_14_1, s_3_15_1; 
    wire s_1_14_1; 
    wire s_2_15_1, s_3_16_1; 
    wire s_1_15_1; 
    wire s_2_16_1, s_3_17_1; 
    wire s_1_16_1; 
    wire s_2_17_1, s_3_18_1; 
    wire s_1_17_1; 
    wire s_2_18_1, s_3_19_1; 
    wire s_1_18_1; 
    wire s_2_19_1, s_3_20_1; 
    wire s_1_19_1; 
    wire s_2_20_1, s_3_21_1; 
    wire s_1_20_1; 
    wire s_2_21_1, s_3_22_1; 
    wire s_1_21_1; 
    wire s_2_22_1, s_3_23_1; 
    wire s_1_22_1; 
    wire s_2_23_1, s_3_24_1; 
    wire s_1_23_1; 
    wire s_2_24_1, s_3_25_1; 
    wire s_1_24_1; 
    wire s_2_25_1, s_3_26_1; 
    wire s_1_25_1; 
    wire s_2_26_1, s_3_27_1; 
    wire s_1_26_1; 
    wire s_2_27_1, s_3_28_1; 
    wire s_1_27_1; 
    wire s_2_28_1, s_3_29_1; 
    wire s_1_28_1; 
    wire s_2_29_1, s_3_30_1; 
    wire s_1_29_1; 
    wire s_2_30_1, s_3_31_1; 
    wire s_1_30_1; 
    wire s_2_31_1, s_3_32_1; 
    wire s_1_31_1; 
    wire s_2_32_1, s_3_33_1; 
    wire s_1_32_1; 
    // total 1 half adders and 28 full adders
    // d_2 = 3 done

    wire s_1_1_0, s_2_2_0, s_1_2_0; 
    wire s_2_3_0, s_2_4_0; 
    wire s_1_3_0; 
    wire s_1_4_0, s_2_5_0; 
    wire s_1_5_0, s_2_6_0; 
    wire s_1_6_0, s_2_7_0; 
    wire s_1_7_0, s_2_8_0; 
    wire s_1_8_0, s_2_9_0; 
    wire s_1_9_0, s_2_10_0; 
    wire s_1_10_0, s_2_11_0; 
    wire s_1_11_0, s_2_12_0; 
    wire s_1_12_0, s_2_13_0; 
    wire s_1_13_0, s_2_14_0; 
    wire s_1_14_0, s_2_15_0; 
    wire s_1_15_0, s_2_16_0; 
    wire s_1_16_0, s_2_17_0; 
    wire s_1_17_0, s_2_18_0; 
    wire s_1_18_0, s_2_19_0; 
    wire s_1_19_0, s_2_20_0; 
    wire s_1_20_0, s_2_21_0; 
    wire s_1_21_0, s_2_22_0; 
    wire s_1_22_0, s_2_23_0; 
    wire s_1_23_0, s_2_24_0; 
    wire s_1_24_0, s_2_25_0; 
    wire s_1_25_0, s_2_26_0; 
    wire s_1_26_0, s_2_27_0; 
    wire s_1_27_0, s_2_28_0; 
    wire s_1_28_0, s_2_29_0; 
    wire s_1_29_0, s_2_30_0; 
    wire s_1_30_0, s_2_31_0; 
    wire s_1_31_0, s_2_32_0; 
    wire s_1_32_0, s_2_33_0; 
    // total 1 half adders and 29 full adders
    // d_1 = 2 done

    assign s_1_1_8 = A[0] & B[0];
    assign s_1_2_8 = A[0] & B[1];
    assign s_1_3_8 = A[0] & B[2];
    assign s_1_4_8 = A[0] & B[3];
    assign s_1_5_8 = A[0] & B[4];
    assign s_1_6_8 = A[0] & B[5];
    assign s_1_7_8 = A[0] & B[6];
    assign s_1_8_8 = A[0] & B[7];
    assign s_1_9_8 = A[0] & B[8];
    assign s_1_10_8 = A[0] & B[9];
    assign s_1_11_8 = A[0] & B[10];
    assign s_1_12_8 = A[0] & B[11];
    assign s_1_13_8 = A[0] & B[12];
    assign s_1_14_8 = A[0] & B[13];
    assign s_1_15_8 = A[0] & B[14];
    assign s_1_16_8 = A[0] & B[15];
    assign s_1_17_8 = A[0] & B[16];
    assign s_1_18_8 = A[0] & B[17];
    assign s_1_19_8 = A[0] & B[18];
    assign s_1_20_8 = A[0] & B[19];
    assign s_1_21_8 = A[0] & B[20];
    assign s_1_22_8 = A[0] & B[21];
    assign s_1_23_8 = A[0] & B[22];
    assign s_1_24_8 = A[0] & B[23];
    assign s_1_25_8 = A[0] & B[24];
    assign s_1_26_8 = A[0] & B[25];
    assign s_1_27_8 = A[0] & B[26];
    assign s_1_28_8 = A[0] & B[27];
    assign s_1_29_8 = A[0] & B[28];
    assign s_1_30_8 = A[0] & B[29];
    assign s_1_31_8 = A[0] & B[30];
    assign s_1_32_8 = A[0] & B[31];
    assign s_2_2_8 = A[1] & B[0];
    assign s_2_3_8 = A[1] & B[1];
    assign s_2_4_8 = A[1] & B[2];
    assign s_2_5_8 = A[1] & B[3];
    assign s_2_6_8 = A[1] & B[4];
    assign s_2_7_8 = A[1] & B[5];
    assign s_2_8_8 = A[1] & B[6];
    assign s_2_9_8 = A[1] & B[7];
    assign s_2_10_8 = A[1] & B[8];
    assign s_2_11_8 = A[1] & B[9];
    assign s_2_12_8 = A[1] & B[10];
    assign s_2_13_8 = A[1] & B[11];
    assign s_2_14_8 = A[1] & B[12];
    assign s_2_15_8 = A[1] & B[13];
    assign s_2_16_8 = A[1] & B[14];
    assign s_2_17_8 = A[1] & B[15];
    assign s_2_18_8 = A[1] & B[16];
    assign s_2_19_8 = A[1] & B[17];
    assign s_2_20_8 = A[1] & B[18];
    assign s_2_21_8 = A[1] & B[19];
    assign s_2_22_8 = A[1] & B[20];
    assign s_2_23_8 = A[1] & B[21];
    assign s_2_24_8 = A[1] & B[22];
    assign s_2_25_8 = A[1] & B[23];
    assign s_2_26_8 = A[1] & B[24];
    assign s_2_27_8 = A[1] & B[25];
    assign s_2_28_8 = A[1] & B[26];
    assign s_2_29_8 = A[1] & B[27];
    assign s_2_30_8 = A[1] & B[28];
    assign s_2_31_8 = A[1] & B[29];
    assign s_2_32_8 = A[1] & B[30];
    assign s_3_3_8 = A[2] & B[0];
    assign s_3_4_8 = A[2] & B[1];
    assign s_3_5_8 = A[2] & B[2];
    assign s_3_6_8 = A[2] & B[3];
    assign s_3_7_8 = A[2] & B[4];
    assign s_3_8_8 = A[2] & B[5];
    assign s_3_9_8 = A[2] & B[6];
    assign s_3_10_8 = A[2] & B[7];
    assign s_3_11_8 = A[2] & B[8];
    assign s_3_12_8 = A[2] & B[9];
    assign s_3_13_8 = A[2] & B[10];
    assign s_3_14_8 = A[2] & B[11];
    assign s_3_15_8 = A[2] & B[12];
    assign s_3_16_8 = A[2] & B[13];
    assign s_3_17_8 = A[2] & B[14];
    assign s_3_18_8 = A[2] & B[15];
    assign s_3_19_8 = A[2] & B[16];
    assign s_3_20_8 = A[2] & B[17];
    assign s_3_21_8 = A[2] & B[18];
    assign s_3_22_8 = A[2] & B[19];
    assign s_3_23_8 = A[2] & B[20];
    assign s_3_24_8 = A[2] & B[21];
    assign s_3_25_8 = A[2] & B[22];
    assign s_3_26_8 = A[2] & B[23];
    assign s_3_27_8 = A[2] & B[24];
    assign s_3_28_8 = A[2] & B[25];
    assign s_3_29_8 = A[2] & B[26];
    assign s_3_30_8 = A[2] & B[27];
    assign s_3_31_8 = A[2] & B[28];
    assign s_3_32_8 = A[2] & B[29];
    assign s_4_4_8 = A[3] & B[0];
    assign s_4_5_8 = A[3] & B[1];
    assign s_4_6_8 = A[3] & B[2];
    assign s_4_7_8 = A[3] & B[3];
    assign s_4_8_8 = A[3] & B[4];
    assign s_4_9_8 = A[3] & B[5];
    assign s_4_10_8 = A[3] & B[6];
    assign s_4_11_8 = A[3] & B[7];
    assign s_4_12_8 = A[3] & B[8];
    assign s_4_13_8 = A[3] & B[9];
    assign s_4_14_8 = A[3] & B[10];
    assign s_4_15_8 = A[3] & B[11];
    assign s_4_16_8 = A[3] & B[12];
    assign s_4_17_8 = A[3] & B[13];
    assign s_4_18_8 = A[3] & B[14];
    assign s_4_19_8 = A[3] & B[15];
    assign s_4_20_8 = A[3] & B[16];
    assign s_4_21_8 = A[3] & B[17];
    assign s_4_22_8 = A[3] & B[18];
    assign s_4_23_8 = A[3] & B[19];
    assign s_4_24_8 = A[3] & B[20];
    assign s_4_25_8 = A[3] & B[21];
    assign s_4_26_8 = A[3] & B[22];
    assign s_4_27_8 = A[3] & B[23];
    assign s_4_28_8 = A[3] & B[24];
    assign s_4_29_8 = A[3] & B[25];
    assign s_4_30_8 = A[3] & B[26];
    assign s_4_31_8 = A[3] & B[27];
    assign s_4_32_8 = A[3] & B[28];
    assign s_5_5_8 = A[4] & B[0];
    assign s_5_6_8 = A[4] & B[1];
    assign s_5_7_8 = A[4] & B[2];
    assign s_5_8_8 = A[4] & B[3];
    assign s_5_9_8 = A[4] & B[4];
    assign s_5_10_8 = A[4] & B[5];
    assign s_5_11_8 = A[4] & B[6];
    assign s_5_12_8 = A[4] & B[7];
    assign s_5_13_8 = A[4] & B[8];
    assign s_5_14_8 = A[4] & B[9];
    assign s_5_15_8 = A[4] & B[10];
    assign s_5_16_8 = A[4] & B[11];
    assign s_5_17_8 = A[4] & B[12];
    assign s_5_18_8 = A[4] & B[13];
    assign s_5_19_8 = A[4] & B[14];
    assign s_5_20_8 = A[4] & B[15];
    assign s_5_21_8 = A[4] & B[16];
    assign s_5_22_8 = A[4] & B[17];
    assign s_5_23_8 = A[4] & B[18];
    assign s_5_24_8 = A[4] & B[19];
    assign s_5_25_8 = A[4] & B[20];
    assign s_5_26_8 = A[4] & B[21];
    assign s_5_27_8 = A[4] & B[22];
    assign s_5_28_8 = A[4] & B[23];
    assign s_5_29_8 = A[4] & B[24];
    assign s_5_30_8 = A[4] & B[25];
    assign s_5_31_8 = A[4] & B[26];
    assign s_5_32_8 = A[4] & B[27];
    assign s_6_6_8 = A[5] & B[0];
    assign s_6_7_8 = A[5] & B[1];
    assign s_6_8_8 = A[5] & B[2];
    assign s_6_9_8 = A[5] & B[3];
    assign s_6_10_8 = A[5] & B[4];
    assign s_6_11_8 = A[5] & B[5];
    assign s_6_12_8 = A[5] & B[6];
    assign s_6_13_8 = A[5] & B[7];
    assign s_6_14_8 = A[5] & B[8];
    assign s_6_15_8 = A[5] & B[9];
    assign s_6_16_8 = A[5] & B[10];
    assign s_6_17_8 = A[5] & B[11];
    assign s_6_18_8 = A[5] & B[12];
    assign s_6_19_8 = A[5] & B[13];
    assign s_6_20_8 = A[5] & B[14];
    assign s_6_21_8 = A[5] & B[15];
    assign s_6_22_8 = A[5] & B[16];
    assign s_6_23_8 = A[5] & B[17];
    assign s_6_24_8 = A[5] & B[18];
    assign s_6_25_8 = A[5] & B[19];
    assign s_6_26_8 = A[5] & B[20];
    assign s_6_27_8 = A[5] & B[21];
    assign s_6_28_8 = A[5] & B[22];
    assign s_6_29_8 = A[5] & B[23];
    assign s_6_30_8 = A[5] & B[24];
    assign s_6_31_8 = A[5] & B[25];
    assign s_6_32_8 = A[5] & B[26];
    assign s_7_7_8 = A[6] & B[0];
    assign s_7_8_8 = A[6] & B[1];
    assign s_7_9_8 = A[6] & B[2];
    assign s_7_10_8 = A[6] & B[3];
    assign s_7_11_8 = A[6] & B[4];
    assign s_7_12_8 = A[6] & B[5];
    assign s_7_13_8 = A[6] & B[6];
    assign s_7_14_8 = A[6] & B[7];
    assign s_7_15_8 = A[6] & B[8];
    assign s_7_16_8 = A[6] & B[9];
    assign s_7_17_8 = A[6] & B[10];
    assign s_7_18_8 = A[6] & B[11];
    assign s_7_19_8 = A[6] & B[12];
    assign s_7_20_8 = A[6] & B[13];
    assign s_7_21_8 = A[6] & B[14];
    assign s_7_22_8 = A[6] & B[15];
    assign s_7_23_8 = A[6] & B[16];
    assign s_7_24_8 = A[6] & B[17];
    assign s_7_25_8 = A[6] & B[18];
    assign s_7_26_8 = A[6] & B[19];
    assign s_7_27_8 = A[6] & B[20];
    assign s_7_28_8 = A[6] & B[21];
    assign s_7_29_8 = A[6] & B[22];
    assign s_7_30_8 = A[6] & B[23];
    assign s_7_31_8 = A[6] & B[24];
    assign s_7_32_8 = A[6] & B[25];
    assign s_8_8_8 = A[7] & B[0];
    assign s_8_9_8 = A[7] & B[1];
    assign s_8_10_8 = A[7] & B[2];
    assign s_8_11_8 = A[7] & B[3];
    assign s_8_12_8 = A[7] & B[4];
    assign s_8_13_8 = A[7] & B[5];
    assign s_8_14_8 = A[7] & B[6];
    assign s_8_15_8 = A[7] & B[7];
    assign s_8_16_8 = A[7] & B[8];
    assign s_8_17_8 = A[7] & B[9];
    assign s_8_18_8 = A[7] & B[10];
    assign s_8_19_8 = A[7] & B[11];
    assign s_8_20_8 = A[7] & B[12];
    assign s_8_21_8 = A[7] & B[13];
    assign s_8_22_8 = A[7] & B[14];
    assign s_8_23_8 = A[7] & B[15];
    assign s_8_24_8 = A[7] & B[16];
    assign s_8_25_8 = A[7] & B[17];
    assign s_8_26_8 = A[7] & B[18];
    assign s_8_27_8 = A[7] & B[19];
    assign s_8_28_8 = A[7] & B[20];
    assign s_8_29_8 = A[7] & B[21];
    assign s_8_30_8 = A[7] & B[22];
    assign s_8_31_8 = A[7] & B[23];
    assign s_8_32_8 = A[7] & B[24];
    assign s_9_9_8 = A[8] & B[0];
    assign s_9_10_8 = A[8] & B[1];
    assign s_9_11_8 = A[8] & B[2];
    assign s_9_12_8 = A[8] & B[3];
    assign s_9_13_8 = A[8] & B[4];
    assign s_9_14_8 = A[8] & B[5];
    assign s_9_15_8 = A[8] & B[6];
    assign s_9_16_8 = A[8] & B[7];
    assign s_9_17_8 = A[8] & B[8];
    assign s_9_18_8 = A[8] & B[9];
    assign s_9_19_8 = A[8] & B[10];
    assign s_9_20_8 = A[8] & B[11];
    assign s_9_21_8 = A[8] & B[12];
    assign s_9_22_8 = A[8] & B[13];
    assign s_9_23_8 = A[8] & B[14];
    assign s_9_24_8 = A[8] & B[15];
    assign s_9_25_8 = A[8] & B[16];
    assign s_9_26_8 = A[8] & B[17];
    assign s_9_27_8 = A[8] & B[18];
    assign s_9_28_8 = A[8] & B[19];
    assign s_9_29_8 = A[8] & B[20];
    assign s_9_30_8 = A[8] & B[21];
    assign s_9_31_8 = A[8] & B[22];
    assign s_9_32_8 = A[8] & B[23];
    assign s_10_10_8 = A[9] & B[0];
    assign s_10_11_8 = A[9] & B[1];
    assign s_10_12_8 = A[9] & B[2];
    assign s_10_13_8 = A[9] & B[3];
    assign s_10_14_8 = A[9] & B[4];
    assign s_10_15_8 = A[9] & B[5];
    assign s_10_16_8 = A[9] & B[6];
    assign s_10_17_8 = A[9] & B[7];
    assign s_10_18_8 = A[9] & B[8];
    assign s_10_19_8 = A[9] & B[9];
    assign s_10_20_8 = A[9] & B[10];
    assign s_10_21_8 = A[9] & B[11];
    assign s_10_22_8 = A[9] & B[12];
    assign s_10_23_8 = A[9] & B[13];
    assign s_10_24_8 = A[9] & B[14];
    assign s_10_25_8 = A[9] & B[15];
    assign s_10_26_8 = A[9] & B[16];
    assign s_10_27_8 = A[9] & B[17];
    assign s_10_28_8 = A[9] & B[18];
    assign s_10_29_8 = A[9] & B[19];
    assign s_10_30_8 = A[9] & B[20];
    assign s_10_31_8 = A[9] & B[21];
    assign s_10_32_8 = A[9] & B[22];
    assign s_11_11_8 = A[10] & B[0];
    assign s_11_12_8 = A[10] & B[1];
    assign s_11_13_8 = A[10] & B[2];
    assign s_11_14_8 = A[10] & B[3];
    assign s_11_15_8 = A[10] & B[4];
    assign s_11_16_8 = A[10] & B[5];
    assign s_11_17_8 = A[10] & B[6];
    assign s_11_18_8 = A[10] & B[7];
    assign s_11_19_8 = A[10] & B[8];
    assign s_11_20_8 = A[10] & B[9];
    assign s_11_21_8 = A[10] & B[10];
    assign s_11_22_8 = A[10] & B[11];
    assign s_11_23_8 = A[10] & B[12];
    assign s_11_24_8 = A[10] & B[13];
    assign s_11_25_8 = A[10] & B[14];
    assign s_11_26_8 = A[10] & B[15];
    assign s_11_27_8 = A[10] & B[16];
    assign s_11_28_8 = A[10] & B[17];
    assign s_11_29_8 = A[10] & B[18];
    assign s_11_30_8 = A[10] & B[19];
    assign s_11_31_8 = A[10] & B[20];
    assign s_11_32_8 = A[10] & B[21];
    assign s_12_12_8 = A[11] & B[0];
    assign s_12_13_8 = A[11] & B[1];
    assign s_12_14_8 = A[11] & B[2];
    assign s_12_15_8 = A[11] & B[3];
    assign s_12_16_8 = A[11] & B[4];
    assign s_12_17_8 = A[11] & B[5];
    assign s_12_18_8 = A[11] & B[6];
    assign s_12_19_8 = A[11] & B[7];
    assign s_12_20_8 = A[11] & B[8];
    assign s_12_21_8 = A[11] & B[9];
    assign s_12_22_8 = A[11] & B[10];
    assign s_12_23_8 = A[11] & B[11];
    assign s_12_24_8 = A[11] & B[12];
    assign s_12_25_8 = A[11] & B[13];
    assign s_12_26_8 = A[11] & B[14];
    assign s_12_27_8 = A[11] & B[15];
    assign s_12_28_8 = A[11] & B[16];
    assign s_12_29_8 = A[11] & B[17];
    assign s_12_30_8 = A[11] & B[18];
    assign s_12_31_8 = A[11] & B[19];
    assign s_12_32_8 = A[11] & B[20];
    assign s_13_13_8 = A[12] & B[0];
    assign s_13_14_8 = A[12] & B[1];
    assign s_13_15_8 = A[12] & B[2];
    assign s_13_16_8 = A[12] & B[3];
    assign s_13_17_8 = A[12] & B[4];
    assign s_13_18_8 = A[12] & B[5];
    assign s_13_19_8 = A[12] & B[6];
    assign s_13_20_8 = A[12] & B[7];
    assign s_13_21_8 = A[12] & B[8];
    assign s_13_22_8 = A[12] & B[9];
    assign s_13_23_8 = A[12] & B[10];
    assign s_13_24_8 = A[12] & B[11];
    assign s_13_25_8 = A[12] & B[12];
    assign s_13_26_8 = A[12] & B[13];
    assign s_13_27_8 = A[12] & B[14];
    assign s_13_28_8 = A[12] & B[15];
    assign s_13_29_8 = A[12] & B[16];
    assign s_13_30_8 = A[12] & B[17];
    assign s_13_31_8 = A[12] & B[18];
    assign s_13_32_8 = A[12] & B[19];
    assign s_14_14_8 = A[13] & B[0];
    assign s_14_15_8 = A[13] & B[1];
    assign s_14_16_8 = A[13] & B[2];
    assign s_14_17_8 = A[13] & B[3];
    assign s_14_18_8 = A[13] & B[4];
    assign s_14_19_8 = A[13] & B[5];
    assign s_14_20_8 = A[13] & B[6];
    assign s_14_21_8 = A[13] & B[7];
    assign s_14_22_8 = A[13] & B[8];
    assign s_14_23_8 = A[13] & B[9];
    assign s_14_24_8 = A[13] & B[10];
    assign s_14_25_8 = A[13] & B[11];
    assign s_14_26_8 = A[13] & B[12];
    assign s_14_27_8 = A[13] & B[13];
    assign s_14_28_8 = A[13] & B[14];
    assign s_14_29_8 = A[13] & B[15];
    assign s_14_30_8 = A[13] & B[16];
    assign s_14_31_8 = A[13] & B[17];
    assign s_14_32_8 = A[13] & B[18];
    assign s_15_15_8 = A[14] & B[0];
    assign s_15_16_8 = A[14] & B[1];
    assign s_15_17_8 = A[14] & B[2];
    assign s_15_18_8 = A[14] & B[3];
    assign s_15_19_8 = A[14] & B[4];
    assign s_15_20_8 = A[14] & B[5];
    assign s_15_21_8 = A[14] & B[6];
    assign s_15_22_8 = A[14] & B[7];
    assign s_15_23_8 = A[14] & B[8];
    assign s_15_24_8 = A[14] & B[9];
    assign s_15_25_8 = A[14] & B[10];
    assign s_15_26_8 = A[14] & B[11];
    assign s_15_27_8 = A[14] & B[12];
    assign s_15_28_8 = A[14] & B[13];
    assign s_15_29_8 = A[14] & B[14];
    assign s_15_30_8 = A[14] & B[15];
    assign s_15_31_8 = A[14] & B[16];
    assign s_15_32_8 = A[14] & B[17];
    assign s_16_16_8 = A[15] & B[0];
    assign s_16_17_8 = A[15] & B[1];
    assign s_16_18_8 = A[15] & B[2];
    assign s_16_19_8 = A[15] & B[3];
    assign s_16_20_8 = A[15] & B[4];
    assign s_16_21_8 = A[15] & B[5];
    assign s_16_22_8 = A[15] & B[6];
    assign s_16_23_8 = A[15] & B[7];
    assign s_16_24_8 = A[15] & B[8];
    assign s_16_25_8 = A[15] & B[9];
    assign s_16_26_8 = A[15] & B[10];
    assign s_16_27_8 = A[15] & B[11];
    assign s_16_28_8 = A[15] & B[12];
    assign s_16_29_8 = A[15] & B[13];
    assign s_16_30_8 = A[15] & B[14];
    assign s_16_31_8 = A[15] & B[15];
    assign s_16_32_8 = A[15] & B[16];
    assign s_17_17_8 = A[16] & B[0];
    assign s_17_18_8 = A[16] & B[1];
    assign s_17_19_8 = A[16] & B[2];
    assign s_17_20_8 = A[16] & B[3];
    assign s_17_21_8 = A[16] & B[4];
    assign s_17_22_8 = A[16] & B[5];
    assign s_17_23_8 = A[16] & B[6];
    assign s_17_24_8 = A[16] & B[7];
    assign s_17_25_8 = A[16] & B[8];
    assign s_17_26_8 = A[16] & B[9];
    assign s_17_27_8 = A[16] & B[10];
    assign s_17_28_8 = A[16] & B[11];
    assign s_17_29_8 = A[16] & B[12];
    assign s_17_30_8 = A[16] & B[13];
    assign s_17_31_8 = A[16] & B[14];
    assign s_17_32_8 = A[16] & B[15];
    assign s_18_18_8 = A[17] & B[0];
    assign s_18_19_8 = A[17] & B[1];
    assign s_18_20_8 = A[17] & B[2];
    assign s_18_21_8 = A[17] & B[3];
    assign s_18_22_8 = A[17] & B[4];
    assign s_18_23_8 = A[17] & B[5];
    assign s_18_24_8 = A[17] & B[6];
    assign s_18_25_8 = A[17] & B[7];
    assign s_18_26_8 = A[17] & B[8];
    assign s_18_27_8 = A[17] & B[9];
    assign s_18_28_8 = A[17] & B[10];
    assign s_18_29_8 = A[17] & B[11];
    assign s_18_30_8 = A[17] & B[12];
    assign s_18_31_8 = A[17] & B[13];
    assign s_18_32_8 = A[17] & B[14];
    assign s_19_19_8 = A[18] & B[0];
    assign s_19_20_8 = A[18] & B[1];
    assign s_19_21_8 = A[18] & B[2];
    assign s_19_22_8 = A[18] & B[3];
    assign s_19_23_8 = A[18] & B[4];
    assign s_19_24_8 = A[18] & B[5];
    assign s_19_25_8 = A[18] & B[6];
    assign s_19_26_8 = A[18] & B[7];
    assign s_19_27_8 = A[18] & B[8];
    assign s_19_28_8 = A[18] & B[9];
    assign s_19_29_8 = A[18] & B[10];
    assign s_19_30_8 = A[18] & B[11];
    assign s_19_31_8 = A[18] & B[12];
    assign s_19_32_8 = A[18] & B[13];
    assign s_20_20_8 = A[19] & B[0];
    assign s_20_21_8 = A[19] & B[1];
    assign s_20_22_8 = A[19] & B[2];
    assign s_20_23_8 = A[19] & B[3];
    assign s_20_24_8 = A[19] & B[4];
    assign s_20_25_8 = A[19] & B[5];
    assign s_20_26_8 = A[19] & B[6];
    assign s_20_27_8 = A[19] & B[7];
    assign s_20_28_8 = A[19] & B[8];
    assign s_20_29_8 = A[19] & B[9];
    assign s_20_30_8 = A[19] & B[10];
    assign s_20_31_8 = A[19] & B[11];
    assign s_20_32_8 = A[19] & B[12];
    assign s_21_21_8 = A[20] & B[0];
    assign s_21_22_8 = A[20] & B[1];
    assign s_21_23_8 = A[20] & B[2];
    assign s_21_24_8 = A[20] & B[3];
    assign s_21_25_8 = A[20] & B[4];
    assign s_21_26_8 = A[20] & B[5];
    assign s_21_27_8 = A[20] & B[6];
    assign s_21_28_8 = A[20] & B[7];
    assign s_21_29_8 = A[20] & B[8];
    assign s_21_30_8 = A[20] & B[9];
    assign s_21_31_8 = A[20] & B[10];
    assign s_21_32_8 = A[20] & B[11];
    assign s_22_22_8 = A[21] & B[0];
    assign s_22_23_8 = A[21] & B[1];
    assign s_22_24_8 = A[21] & B[2];
    assign s_22_25_8 = A[21] & B[3];
    assign s_22_26_8 = A[21] & B[4];
    assign s_22_27_8 = A[21] & B[5];
    assign s_22_28_8 = A[21] & B[6];
    assign s_22_29_8 = A[21] & B[7];
    assign s_22_30_8 = A[21] & B[8];
    assign s_22_31_8 = A[21] & B[9];
    assign s_22_32_8 = A[21] & B[10];
    assign s_23_23_8 = A[22] & B[0];
    assign s_23_24_8 = A[22] & B[1];
    assign s_23_25_8 = A[22] & B[2];
    assign s_23_26_8 = A[22] & B[3];
    assign s_23_27_8 = A[22] & B[4];
    assign s_23_28_8 = A[22] & B[5];
    assign s_23_29_8 = A[22] & B[6];
    assign s_23_30_8 = A[22] & B[7];
    assign s_23_31_8 = A[22] & B[8];
    assign s_23_32_8 = A[22] & B[9];
    assign s_24_24_8 = A[23] & B[0];
    assign s_24_25_8 = A[23] & B[1];
    assign s_24_26_8 = A[23] & B[2];
    assign s_24_27_8 = A[23] & B[3];
    assign s_24_28_8 = A[23] & B[4];
    assign s_24_29_8 = A[23] & B[5];
    assign s_24_30_8 = A[23] & B[6];
    assign s_24_31_8 = A[23] & B[7];
    assign s_24_32_8 = A[23] & B[8];
    assign s_25_25_8 = A[24] & B[0];
    assign s_25_26_8 = A[24] & B[1];
    assign s_25_27_8 = A[24] & B[2];
    assign s_25_28_8 = A[24] & B[3];
    assign s_25_29_8 = A[24] & B[4];
    assign s_25_30_8 = A[24] & B[5];
    assign s_25_31_8 = A[24] & B[6];
    assign s_25_32_8 = A[24] & B[7];
    assign s_26_26_8 = A[25] & B[0];
    assign s_26_27_8 = A[25] & B[1];
    assign s_26_28_8 = A[25] & B[2];
    assign s_26_29_8 = A[25] & B[3];
    assign s_26_30_8 = A[25] & B[4];
    assign s_26_31_8 = A[25] & B[5];
    assign s_26_32_8 = A[25] & B[6];
    assign s_27_27_8 = A[26] & B[0];
    assign s_27_28_8 = A[26] & B[1];
    assign s_27_29_8 = A[26] & B[2];
    assign s_27_30_8 = A[26] & B[3];
    assign s_27_31_8 = A[26] & B[4];
    assign s_27_32_8 = A[26] & B[5];
    assign s_28_28_8 = A[27] & B[0];
    assign s_28_29_8 = A[27] & B[1];
    assign s_28_30_8 = A[27] & B[2];
    assign s_28_31_8 = A[27] & B[3];
    assign s_28_32_8 = A[27] & B[4];
    assign s_29_29_8 = A[28] & B[0];
    assign s_29_30_8 = A[28] & B[1];
    assign s_29_31_8 = A[28] & B[2];
    assign s_29_32_8 = A[28] & B[3];
    assign s_30_30_8 = A[29] & B[0];
    assign s_30_31_8 = A[29] & B[1];
    assign s_30_32_8 = A[29] & B[2];
    assign s_31_31_8 = A[30] & B[0];
    assign s_31_32_8 = A[30] & B[1];
    assign s_32_32_8 = A[31] & B[0];

    assign s_1_1_7 = s_1_1_8;
    assign s_2_2_7 = s_1_2_8;
    assign s_1_2_7 = s_2_2_8;
    assign s_3_3_7 = s_1_3_8;
    assign s_2_3_7 = s_2_3_8;
    assign s_1_3_7 = s_3_3_8;
    assign s_4_4_7 = s_1_4_8;
    assign s_3_4_7 = s_2_4_8;
    assign s_2_4_7 = s_3_4_8;
    assign s_1_4_7 = s_4_4_8;
    assign s_5_5_7 = s_1_5_8;
    assign s_4_5_7 = s_2_5_8;
    assign s_3_5_7 = s_3_5_8;
    assign s_2_5_7 = s_4_5_8;
    assign s_1_5_7 = s_5_5_8;
    assign s_6_6_7 = s_1_6_8;
    assign s_5_6_7 = s_2_6_8;
    assign s_4_6_7 = s_3_6_8;
    assign s_3_6_7 = s_4_6_8;
    assign s_2_6_7 = s_5_6_8;
    assign s_1_6_7 = s_6_6_8;
    assign s_7_7_7 = s_1_7_8;
    assign s_6_7_7 = s_2_7_8;
    assign s_5_7_7 = s_3_7_8;
    assign s_4_7_7 = s_4_7_8;
    assign s_3_7_7 = s_5_7_8;
    assign s_2_7_7 = s_6_7_8;
    assign s_1_7_7 = s_7_7_8;
    assign s_8_8_7 = s_1_8_8;
    assign s_7_8_7 = s_2_8_8;
    assign s_6_8_7 = s_3_8_8;
    assign s_5_8_7 = s_4_8_8;
    assign s_4_8_7 = s_5_8_8;
    assign s_3_8_7 = s_6_8_8;
    assign s_2_8_7 = s_7_8_8;
    assign s_1_8_7 = s_8_8_8;
    assign s_9_9_7 = s_1_9_8;
    assign s_8_9_7 = s_2_9_8;
    assign s_7_9_7 = s_3_9_8;
    assign s_6_9_7 = s_4_9_8;
    assign s_5_9_7 = s_5_9_8;
    assign s_4_9_7 = s_6_9_8;
    assign s_3_9_7 = s_7_9_8;
    assign s_2_9_7 = s_8_9_8;
    assign s_1_9_7 = s_9_9_8;
    assign s_10_10_7 = s_1_10_8;
    assign s_9_10_7 = s_2_10_8;
    assign s_8_10_7 = s_3_10_8;
    assign s_7_10_7 = s_4_10_8;
    assign s_6_10_7 = s_5_10_8;
    assign s_5_10_7 = s_6_10_8;
    assign s_4_10_7 = s_7_10_8;
    assign s_3_10_7 = s_8_10_8;
    assign s_2_10_7 = s_9_10_8;
    assign s_1_10_7 = s_10_10_8;
    assign s_11_11_7 = s_1_11_8;
    assign s_10_11_7 = s_2_11_8;
    assign s_9_11_7 = s_3_11_8;
    assign s_8_11_7 = s_4_11_8;
    assign s_7_11_7 = s_5_11_8;
    assign s_6_11_7 = s_6_11_8;
    assign s_5_11_7 = s_7_11_8;
    assign s_4_11_7 = s_8_11_8;
    assign s_3_11_7 = s_9_11_8;
    assign s_2_11_7 = s_10_11_8;
    assign s_1_11_7 = s_11_11_8;
    assign s_12_12_7 = s_1_12_8;
    assign s_11_12_7 = s_2_12_8;
    assign s_10_12_7 = s_3_12_8;
    assign s_9_12_7 = s_4_12_8;
    assign s_8_12_7 = s_5_12_8;
    assign s_7_12_7 = s_6_12_8;
    assign s_6_12_7 = s_7_12_8;
    assign s_5_12_7 = s_8_12_8;
    assign s_4_12_7 = s_9_12_8;
    assign s_3_12_7 = s_10_12_8;
    assign s_2_12_7 = s_11_12_8;
    assign s_1_12_7 = s_12_12_8;
    assign s_13_13_7 = s_1_13_8;
    assign s_12_13_7 = s_2_13_8;
    assign s_11_13_7 = s_3_13_8;
    assign s_10_13_7 = s_4_13_8;
    assign s_9_13_7 = s_5_13_8;
    assign s_8_13_7 = s_6_13_8;
    assign s_7_13_7 = s_7_13_8;
    assign s_6_13_7 = s_8_13_8;
    assign s_5_13_7 = s_9_13_8;
    assign s_4_13_7 = s_10_13_8;
    assign s_3_13_7 = s_11_13_8;
    assign s_2_13_7 = s_12_13_8;
    assign s_1_13_7 = s_13_13_8;
    assign s_14_14_7 = s_1_14_8;
    assign s_13_14_7 = s_2_14_8;
    assign s_12_14_7 = s_3_14_8;
    assign s_11_14_7 = s_4_14_8;
    assign s_10_14_7 = s_5_14_8;
    assign s_9_14_7 = s_6_14_8;
    assign s_8_14_7 = s_7_14_8;
    assign s_7_14_7 = s_8_14_8;
    assign s_6_14_7 = s_9_14_8;
    assign s_5_14_7 = s_10_14_8;
    assign s_4_14_7 = s_11_14_8;
    assign s_3_14_7 = s_12_14_8;
    assign s_2_14_7 = s_13_14_8;
    assign s_1_14_7 = s_14_14_8;
    assign s_15_15_7 = s_1_15_8;
    assign s_14_15_7 = s_2_15_8;
    assign s_13_15_7 = s_3_15_8;
    assign s_12_15_7 = s_4_15_8;
    assign s_11_15_7 = s_5_15_8;
    assign s_10_15_7 = s_6_15_8;
    assign s_9_15_7 = s_7_15_8;
    assign s_8_15_7 = s_8_15_8;
    assign s_7_15_7 = s_9_15_8;
    assign s_6_15_7 = s_10_15_8;
    assign s_5_15_7 = s_11_15_8;
    assign s_4_15_7 = s_12_15_8;
    assign s_3_15_7 = s_13_15_8;
    assign s_2_15_7 = s_14_15_8;
    assign s_1_15_7 = s_15_15_8;
    assign s_16_16_7 = s_1_16_8;
    assign s_15_16_7 = s_2_16_8;
    assign s_14_16_7 = s_3_16_8;
    assign s_13_16_7 = s_4_16_8;
    assign s_12_16_7 = s_5_16_8;
    assign s_11_16_7 = s_6_16_8;
    assign s_10_16_7 = s_7_16_8;
    assign s_9_16_7 = s_8_16_8;
    assign s_8_16_7 = s_9_16_8;
    assign s_7_16_7 = s_10_16_8;
    assign s_6_16_7 = s_11_16_8;
    assign s_5_16_7 = s_12_16_8;
    assign s_4_16_7 = s_13_16_8;
    assign s_3_16_7 = s_14_16_8;
    assign s_2_16_7 = s_15_16_8;
    assign s_1_16_7 = s_16_16_8;
    assign s_17_17_7 = s_1_17_8;
    assign s_16_17_7 = s_2_17_8;
    assign s_15_17_7 = s_3_17_8;
    assign s_14_17_7 = s_4_17_8;
    assign s_13_17_7 = s_5_17_8;
    assign s_12_17_7 = s_6_17_8;
    assign s_11_17_7 = s_7_17_8;
    assign s_10_17_7 = s_8_17_8;
    assign s_9_17_7 = s_9_17_8;
    assign s_8_17_7 = s_10_17_8;
    assign s_7_17_7 = s_11_17_8;
    assign s_6_17_7 = s_12_17_8;
    assign s_5_17_7 = s_13_17_8;
    assign s_4_17_7 = s_14_17_8;
    assign s_3_17_7 = s_15_17_8;
    assign s_2_17_7 = s_16_17_8;
    assign s_1_17_7 = s_17_17_8;
    assign s_18_18_7 = s_1_18_8;
    assign s_17_18_7 = s_2_18_8;
    assign s_16_18_7 = s_3_18_8;
    assign s_15_18_7 = s_4_18_8;
    assign s_14_18_7 = s_5_18_8;
    assign s_13_18_7 = s_6_18_8;
    assign s_12_18_7 = s_7_18_8;
    assign s_11_18_7 = s_8_18_8;
    assign s_10_18_7 = s_9_18_8;
    assign s_9_18_7 = s_10_18_8;
    assign s_8_18_7 = s_11_18_8;
    assign s_7_18_7 = s_12_18_8;
    assign s_6_18_7 = s_13_18_8;
    assign s_5_18_7 = s_14_18_8;
    assign s_4_18_7 = s_15_18_8;
    assign s_3_18_7 = s_16_18_8;
    assign s_2_18_7 = s_17_18_8;
    assign s_1_18_7 = s_18_18_8;
    assign s_19_19_7 = s_1_19_8;
    assign s_18_19_7 = s_2_19_8;
    assign s_17_19_7 = s_3_19_8;
    assign s_16_19_7 = s_4_19_8;
    assign s_15_19_7 = s_5_19_8;
    assign s_14_19_7 = s_6_19_8;
    assign s_13_19_7 = s_7_19_8;
    assign s_12_19_7 = s_8_19_8;
    assign s_11_19_7 = s_9_19_8;
    assign s_10_19_7 = s_10_19_8;
    assign s_9_19_7 = s_11_19_8;
    assign s_8_19_7 = s_12_19_8;
    assign s_7_19_7 = s_13_19_8;
    assign s_6_19_7 = s_14_19_8;
    assign s_5_19_7 = s_15_19_8;
    assign s_4_19_7 = s_16_19_8;
    assign s_3_19_7 = s_17_19_8;
    assign s_2_19_7 = s_18_19_8;
    assign s_1_19_7 = s_19_19_8;
    assign s_20_20_7 = s_1_20_8;
    assign s_19_20_7 = s_2_20_8;
    assign s_18_20_7 = s_3_20_8;
    assign s_17_20_7 = s_4_20_8;
    assign s_16_20_7 = s_5_20_8;
    assign s_15_20_7 = s_6_20_8;
    assign s_14_20_7 = s_7_20_8;
    assign s_13_20_7 = s_8_20_8;
    assign s_12_20_7 = s_9_20_8;
    assign s_11_20_7 = s_10_20_8;
    assign s_10_20_7 = s_11_20_8;
    assign s_9_20_7 = s_12_20_8;
    assign s_8_20_7 = s_13_20_8;
    assign s_7_20_7 = s_14_20_8;
    assign s_6_20_7 = s_15_20_8;
    assign s_5_20_7 = s_16_20_8;
    assign s_4_20_7 = s_17_20_8;
    assign s_3_20_7 = s_18_20_8;
    assign s_2_20_7 = s_19_20_8;
    assign s_1_20_7 = s_20_20_8;
    assign s_21_21_7 = s_1_21_8;
    assign s_20_21_7 = s_2_21_8;
    assign s_19_21_7 = s_3_21_8;
    assign s_18_21_7 = s_4_21_8;
    assign s_17_21_7 = s_5_21_8;
    assign s_16_21_7 = s_6_21_8;
    assign s_15_21_7 = s_7_21_8;
    assign s_14_21_7 = s_8_21_8;
    assign s_13_21_7 = s_9_21_8;
    assign s_12_21_7 = s_10_21_8;
    assign s_11_21_7 = s_11_21_8;
    assign s_10_21_7 = s_12_21_8;
    assign s_9_21_7 = s_13_21_8;
    assign s_8_21_7 = s_14_21_8;
    assign s_7_21_7 = s_15_21_8;
    assign s_6_21_7 = s_16_21_8;
    assign s_5_21_7 = s_17_21_8;
    assign s_4_21_7 = s_18_21_8;
    assign s_3_21_7 = s_19_21_8;
    assign s_2_21_7 = s_20_21_8;
    assign s_1_21_7 = s_21_21_8;
    assign s_22_22_7 = s_1_22_8;
    assign s_21_22_7 = s_2_22_8;
    assign s_20_22_7 = s_3_22_8;
    assign s_19_22_7 = s_4_22_8;
    assign s_18_22_7 = s_5_22_8;
    assign s_17_22_7 = s_6_22_8;
    assign s_16_22_7 = s_7_22_8;
    assign s_15_22_7 = s_8_22_8;
    assign s_14_22_7 = s_9_22_8;
    assign s_13_22_7 = s_10_22_8;
    assign s_12_22_7 = s_11_22_8;
    assign s_11_22_7 = s_12_22_8;
    assign s_10_22_7 = s_13_22_8;
    assign s_9_22_7 = s_14_22_8;
    assign s_8_22_7 = s_15_22_8;
    assign s_7_22_7 = s_16_22_8;
    assign s_6_22_7 = s_17_22_8;
    assign s_5_22_7 = s_18_22_8;
    assign s_4_22_7 = s_19_22_8;
    assign s_3_22_7 = s_20_22_8;
    assign s_2_22_7 = s_21_22_8;
    assign s_1_22_7 = s_22_22_8;
    assign s_23_23_7 = s_1_23_8;
    assign s_22_23_7 = s_2_23_8;
    assign s_21_23_7 = s_3_23_8;
    assign s_20_23_7 = s_4_23_8;
    assign s_19_23_7 = s_5_23_8;
    assign s_18_23_7 = s_6_23_8;
    assign s_17_23_7 = s_7_23_8;
    assign s_16_23_7 = s_8_23_8;
    assign s_15_23_7 = s_9_23_8;
    assign s_14_23_7 = s_10_23_8;
    assign s_13_23_7 = s_11_23_8;
    assign s_12_23_7 = s_12_23_8;
    assign s_11_23_7 = s_13_23_8;
    assign s_10_23_7 = s_14_23_8;
    assign s_9_23_7 = s_15_23_8;
    assign s_8_23_7 = s_16_23_8;
    assign s_7_23_7 = s_17_23_8;
    assign s_6_23_7 = s_18_23_8;
    assign s_5_23_7 = s_19_23_8;
    assign s_4_23_7 = s_20_23_8;
    assign s_3_23_7 = s_21_23_8;
    assign s_2_23_7 = s_22_23_8;
    assign s_1_23_7 = s_23_23_8;
    assign s_24_24_7 = s_1_24_8;
    assign s_23_24_7 = s_2_24_8;
    assign s_22_24_7 = s_3_24_8;
    assign s_21_24_7 = s_4_24_8;
    assign s_20_24_7 = s_5_24_8;
    assign s_19_24_7 = s_6_24_8;
    assign s_18_24_7 = s_7_24_8;
    assign s_17_24_7 = s_8_24_8;
    assign s_16_24_7 = s_9_24_8;
    assign s_15_24_7 = s_10_24_8;
    assign s_14_24_7 = s_11_24_8;
    assign s_13_24_7 = s_12_24_8;
    assign s_12_24_7 = s_13_24_8;
    assign s_11_24_7 = s_14_24_8;
    assign s_10_24_7 = s_15_24_8;
    assign s_9_24_7 = s_16_24_8;
    assign s_8_24_7 = s_17_24_8;
    assign s_7_24_7 = s_18_24_8;
    assign s_6_24_7 = s_19_24_8;
    assign s_5_24_7 = s_20_24_8;
    assign s_4_24_7 = s_21_24_8;
    assign s_3_24_7 = s_22_24_8;
    assign s_2_24_7 = s_23_24_8;
    assign s_1_24_7 = s_24_24_8;
    assign s_25_25_7 = s_1_25_8;
    assign s_24_25_7 = s_2_25_8;
    assign s_23_25_7 = s_3_25_8;
    assign s_22_25_7 = s_4_25_8;
    assign s_21_25_7 = s_5_25_8;
    assign s_20_25_7 = s_6_25_8;
    assign s_19_25_7 = s_7_25_8;
    assign s_18_25_7 = s_8_25_8;
    assign s_17_25_7 = s_9_25_8;
    assign s_16_25_7 = s_10_25_8;
    assign s_15_25_7 = s_11_25_8;
    assign s_14_25_7 = s_12_25_8;
    assign s_13_25_7 = s_13_25_8;
    assign s_12_25_7 = s_14_25_8;
    assign s_11_25_7 = s_15_25_8;
    assign s_10_25_7 = s_16_25_8;
    assign s_9_25_7 = s_17_25_8;
    assign s_8_25_7 = s_18_25_8;
    assign s_7_25_7 = s_19_25_8;
    assign s_6_25_7 = s_20_25_8;
    assign s_5_25_7 = s_21_25_8;
    assign s_4_25_7 = s_22_25_8;
    assign s_3_25_7 = s_23_25_8;
    assign s_2_25_7 = s_24_25_8;
    assign s_1_25_7 = s_25_25_8;
    assign s_26_26_7 = s_1_26_8;
    assign s_25_26_7 = s_2_26_8;
    assign s_24_26_7 = s_3_26_8;
    assign s_23_26_7 = s_4_26_8;
    assign s_22_26_7 = s_5_26_8;
    assign s_21_26_7 = s_6_26_8;
    assign s_20_26_7 = s_7_26_8;
    assign s_19_26_7 = s_8_26_8;
    assign s_18_26_7 = s_9_26_8;
    assign s_17_26_7 = s_10_26_8;
    assign s_16_26_7 = s_11_26_8;
    assign s_15_26_7 = s_12_26_8;
    assign s_14_26_7 = s_13_26_8;
    assign s_13_26_7 = s_14_26_8;
    assign s_12_26_7 = s_15_26_8;
    assign s_11_26_7 = s_16_26_8;
    assign s_10_26_7 = s_17_26_8;
    assign s_9_26_7 = s_18_26_8;
    assign s_8_26_7 = s_19_26_8;
    assign s_7_26_7 = s_20_26_8;
    assign s_6_26_7 = s_21_26_8;
    assign s_5_26_7 = s_22_26_8;
    assign s_4_26_7 = s_23_26_8;
    assign s_3_26_7 = s_24_26_8;
    assign s_2_26_7 = s_25_26_8;
    assign s_1_26_7 = s_26_26_8;
    assign s_27_27_7 = s_1_27_8;
    assign s_26_27_7 = s_2_27_8;
    assign s_25_27_7 = s_3_27_8;
    assign s_24_27_7 = s_4_27_8;
    assign s_23_27_7 = s_5_27_8;
    assign s_22_27_7 = s_6_27_8;
    assign s_21_27_7 = s_7_27_8;
    assign s_20_27_7 = s_8_27_8;
    assign s_19_27_7 = s_9_27_8;
    assign s_18_27_7 = s_10_27_8;
    assign s_17_27_7 = s_11_27_8;
    assign s_16_27_7 = s_12_27_8;
    assign s_15_27_7 = s_13_27_8;
    assign s_14_27_7 = s_14_27_8;
    assign s_13_27_7 = s_15_27_8;
    assign s_12_27_7 = s_16_27_8;
    assign s_11_27_7 = s_17_27_8;
    assign s_10_27_7 = s_18_27_8;
    assign s_9_27_7 = s_19_27_8;
    assign s_8_27_7 = s_20_27_8;
    assign s_7_27_7 = s_21_27_8;
    assign s_6_27_7 = s_22_27_8;
    assign s_5_27_7 = s_23_27_8;
    assign s_4_27_7 = s_24_27_8;
    assign s_3_27_7 = s_25_27_8;
    assign s_2_27_7 = s_26_27_8;
    assign s_1_27_7 = s_27_27_8;
    assign s_28_28_7 = s_1_28_8;
    assign s_27_28_7 = s_2_28_8;
    assign s_26_28_7 = s_3_28_8;
    assign s_25_28_7 = s_4_28_8;
    assign s_24_28_7 = s_5_28_8;
    assign s_23_28_7 = s_6_28_8;
    assign s_22_28_7 = s_7_28_8;
    assign s_21_28_7 = s_8_28_8;
    assign s_20_28_7 = s_9_28_8;
    assign s_19_28_7 = s_10_28_8;
    assign s_18_28_7 = s_11_28_8;
    assign s_17_28_7 = s_12_28_8;
    assign s_16_28_7 = s_13_28_8;
    assign s_15_28_7 = s_14_28_8;
    assign s_14_28_7 = s_15_28_8;
    assign s_13_28_7 = s_16_28_8;
    assign s_12_28_7 = s_17_28_8;
    assign s_11_28_7 = s_18_28_8;
    assign s_10_28_7 = s_19_28_8;
    assign s_9_28_7 = s_20_28_8;
    assign s_8_28_7 = s_21_28_8;
    assign s_7_28_7 = s_22_28_8;
    assign s_6_28_7 = s_23_28_8;
    assign s_5_28_7 = s_24_28_8;
    assign s_4_28_7 = s_25_28_8;
    assign s_3_28_7 = s_26_28_8;
    assign s_2_28_7 = s_27_28_8;
    assign s_1_28_7 = s_28_28_8;
    HA HA0 (.A(s_1_29_8), .B(s_2_29_8), .S(s_28_29_7), .C(s_28_30_7));
    assign s_27_29_7 = s_3_29_8;
    assign s_26_29_7 = s_4_29_8;
    assign s_25_29_7 = s_5_29_8;
    assign s_24_29_7 = s_6_29_8;
    assign s_23_29_7 = s_7_29_8;
    assign s_22_29_7 = s_8_29_8;
    assign s_21_29_7 = s_9_29_8;
    assign s_20_29_7 = s_10_29_8;
    assign s_19_29_7 = s_11_29_8;
    assign s_18_29_7 = s_12_29_8;
    assign s_17_29_7 = s_13_29_8;
    assign s_16_29_7 = s_14_29_8;
    assign s_15_29_7 = s_15_29_8;
    assign s_14_29_7 = s_16_29_8;
    assign s_13_29_7 = s_17_29_8;
    assign s_12_29_7 = s_18_29_8;
    assign s_11_29_7 = s_19_29_8;
    assign s_10_29_7 = s_20_29_8;
    assign s_9_29_7 = s_21_29_8;
    assign s_8_29_7 = s_22_29_8;
    assign s_7_29_7 = s_23_29_8;
    assign s_6_29_7 = s_24_29_8;
    assign s_5_29_7 = s_25_29_8;
    assign s_4_29_7 = s_26_29_8;
    assign s_3_29_7 = s_27_29_8;
    assign s_2_29_7 = s_28_29_8;
    assign s_1_29_7 = s_29_29_8;
    FA FA0 (.A(s_1_30_8), .B(s_2_30_8), .Cin(s_3_30_8), .S(s_27_30_7), .Cout(s_28_31_7));
    HA HA1 (.A(s_4_30_8), .B(s_5_30_8), .S(s_26_30_7), .C(s_27_31_7));
    assign s_25_30_7 = s_6_30_8;
    assign s_24_30_7 = s_7_30_8;
    assign s_23_30_7 = s_8_30_8;
    assign s_22_30_7 = s_9_30_8;
    assign s_21_30_7 = s_10_30_8;
    assign s_20_30_7 = s_11_30_8;
    assign s_19_30_7 = s_12_30_8;
    assign s_18_30_7 = s_13_30_8;
    assign s_17_30_7 = s_14_30_8;
    assign s_16_30_7 = s_15_30_8;
    assign s_15_30_7 = s_16_30_8;
    assign s_14_30_7 = s_17_30_8;
    assign s_13_30_7 = s_18_30_8;
    assign s_12_30_7 = s_19_30_8;
    assign s_11_30_7 = s_20_30_8;
    assign s_10_30_7 = s_21_30_8;
    assign s_9_30_7 = s_22_30_8;
    assign s_8_30_7 = s_23_30_8;
    assign s_7_30_7 = s_24_30_8;
    assign s_6_30_7 = s_25_30_8;
    assign s_5_30_7 = s_26_30_8;
    assign s_4_30_7 = s_27_30_8;
    assign s_3_30_7 = s_28_30_8;
    assign s_2_30_7 = s_29_30_8;
    assign s_1_30_7 = s_30_30_8;
    FA FA1 (.A(s_1_31_8), .B(s_2_31_8), .Cin(s_3_31_8), .S(s_26_31_7), .Cout(s_28_32_7));
    FA FA2 (.A(s_4_31_8), .B(s_5_31_8), .Cin(s_6_31_8), .S(s_25_31_7), .Cout(s_27_32_7));
    HA HA2 (.A(s_7_31_8), .B(s_8_31_8), .S(s_24_31_7), .C(s_26_32_7));
    assign s_23_31_7 = s_9_31_8;
    assign s_22_31_7 = s_10_31_8;
    assign s_21_31_7 = s_11_31_8;
    assign s_20_31_7 = s_12_31_8;
    assign s_19_31_7 = s_13_31_8;
    assign s_18_31_7 = s_14_31_8;
    assign s_17_31_7 = s_15_31_8;
    assign s_16_31_7 = s_16_31_8;
    assign s_15_31_7 = s_17_31_8;
    assign s_14_31_7 = s_18_31_8;
    assign s_13_31_7 = s_19_31_8;
    assign s_12_31_7 = s_20_31_8;
    assign s_11_31_7 = s_21_31_8;
    assign s_10_31_7 = s_22_31_8;
    assign s_9_31_7 = s_23_31_8;
    assign s_8_31_7 = s_24_31_8;
    assign s_7_31_7 = s_25_31_8;
    assign s_6_31_7 = s_26_31_8;
    assign s_5_31_7 = s_27_31_8;
    assign s_4_31_7 = s_28_31_8;
    assign s_3_31_7 = s_29_31_8;
    assign s_2_31_7 = s_30_31_8;
    assign s_1_31_7 = s_31_31_8;
    FA FA3 (.A(s_1_32_8), .B(s_2_32_8), .Cin(s_3_32_8), .S(s_25_32_7), .Cout(s_28_33_7));
    FA FA4 (.A(s_4_32_8), .B(s_5_32_8), .Cin(s_6_32_8), .S(s_24_32_7), .Cout(s_27_33_7));
    FA FA5 (.A(s_7_32_8), .B(s_8_32_8), .Cin(s_9_32_8), .S(s_23_32_7), .Cout(s_26_33_7));
    HA HA3 (.A(s_10_32_8), .B(s_11_32_8), .S(s_22_32_7), .C(s_25_33_7));
    assign s_21_32_7 = s_12_32_8;
    assign s_20_32_7 = s_13_32_8;
    assign s_19_32_7 = s_14_32_8;
    assign s_18_32_7 = s_15_32_8;
    assign s_17_32_7 = s_16_32_8;
    assign s_16_32_7 = s_17_32_8;
    assign s_15_32_7 = s_18_32_8;
    assign s_14_32_7 = s_19_32_8;
    assign s_13_32_7 = s_20_32_8;
    assign s_12_32_7 = s_21_32_8;
    assign s_11_32_7 = s_22_32_8;
    assign s_10_32_7 = s_23_32_8;
    assign s_9_32_7 = s_24_32_8;
    assign s_8_32_7 = s_25_32_8;
    assign s_7_32_7 = s_26_32_8;
    assign s_6_32_7 = s_27_32_8;
    assign s_5_32_7 = s_28_32_8;
    assign s_4_32_7 = s_29_32_8;
    assign s_3_32_7 = s_30_32_8;
    assign s_2_32_7 = s_31_32_8;
    assign s_1_32_7 = s_32_32_8;
    // total 4 half adders and 6 full adders
    // d_8 = 28 done

    assign s_1_1_6 = s_1_1_7;
    assign s_2_2_6 = s_1_2_7;
    assign s_1_2_6 = s_2_2_7;
    assign s_3_3_6 = s_1_3_7;
    assign s_2_3_6 = s_2_3_7;
    assign s_1_3_6 = s_3_3_7;
    assign s_4_4_6 = s_1_4_7;
    assign s_3_4_6 = s_2_4_7;
    assign s_2_4_6 = s_3_4_7;
    assign s_1_4_6 = s_4_4_7;
    assign s_5_5_6 = s_1_5_7;
    assign s_4_5_6 = s_2_5_7;
    assign s_3_5_6 = s_3_5_7;
    assign s_2_5_6 = s_4_5_7;
    assign s_1_5_6 = s_5_5_7;
    assign s_6_6_6 = s_1_6_7;
    assign s_5_6_6 = s_2_6_7;
    assign s_4_6_6 = s_3_6_7;
    assign s_3_6_6 = s_4_6_7;
    assign s_2_6_6 = s_5_6_7;
    assign s_1_6_6 = s_6_6_7;
    assign s_7_7_6 = s_1_7_7;
    assign s_6_7_6 = s_2_7_7;
    assign s_5_7_6 = s_3_7_7;
    assign s_4_7_6 = s_4_7_7;
    assign s_3_7_6 = s_5_7_7;
    assign s_2_7_6 = s_6_7_7;
    assign s_1_7_6 = s_7_7_7;
    assign s_8_8_6 = s_1_8_7;
    assign s_7_8_6 = s_2_8_7;
    assign s_6_8_6 = s_3_8_7;
    assign s_5_8_6 = s_4_8_7;
    assign s_4_8_6 = s_5_8_7;
    assign s_3_8_6 = s_6_8_7;
    assign s_2_8_6 = s_7_8_7;
    assign s_1_8_6 = s_8_8_7;
    assign s_9_9_6 = s_1_9_7;
    assign s_8_9_6 = s_2_9_7;
    assign s_7_9_6 = s_3_9_7;
    assign s_6_9_6 = s_4_9_7;
    assign s_5_9_6 = s_5_9_7;
    assign s_4_9_6 = s_6_9_7;
    assign s_3_9_6 = s_7_9_7;
    assign s_2_9_6 = s_8_9_7;
    assign s_1_9_6 = s_9_9_7;
    assign s_10_10_6 = s_1_10_7;
    assign s_9_10_6 = s_2_10_7;
    assign s_8_10_6 = s_3_10_7;
    assign s_7_10_6 = s_4_10_7;
    assign s_6_10_6 = s_5_10_7;
    assign s_5_10_6 = s_6_10_7;
    assign s_4_10_6 = s_7_10_7;
    assign s_3_10_6 = s_8_10_7;
    assign s_2_10_6 = s_9_10_7;
    assign s_1_10_6 = s_10_10_7;
    assign s_11_11_6 = s_1_11_7;
    assign s_10_11_6 = s_2_11_7;
    assign s_9_11_6 = s_3_11_7;
    assign s_8_11_6 = s_4_11_7;
    assign s_7_11_6 = s_5_11_7;
    assign s_6_11_6 = s_6_11_7;
    assign s_5_11_6 = s_7_11_7;
    assign s_4_11_6 = s_8_11_7;
    assign s_3_11_6 = s_9_11_7;
    assign s_2_11_6 = s_10_11_7;
    assign s_1_11_6 = s_11_11_7;
    assign s_12_12_6 = s_1_12_7;
    assign s_11_12_6 = s_2_12_7;
    assign s_10_12_6 = s_3_12_7;
    assign s_9_12_6 = s_4_12_7;
    assign s_8_12_6 = s_5_12_7;
    assign s_7_12_6 = s_6_12_7;
    assign s_6_12_6 = s_7_12_7;
    assign s_5_12_6 = s_8_12_7;
    assign s_4_12_6 = s_9_12_7;
    assign s_3_12_6 = s_10_12_7;
    assign s_2_12_6 = s_11_12_7;
    assign s_1_12_6 = s_12_12_7;
    assign s_13_13_6 = s_1_13_7;
    assign s_12_13_6 = s_2_13_7;
    assign s_11_13_6 = s_3_13_7;
    assign s_10_13_6 = s_4_13_7;
    assign s_9_13_6 = s_5_13_7;
    assign s_8_13_6 = s_6_13_7;
    assign s_7_13_6 = s_7_13_7;
    assign s_6_13_6 = s_8_13_7;
    assign s_5_13_6 = s_9_13_7;
    assign s_4_13_6 = s_10_13_7;
    assign s_3_13_6 = s_11_13_7;
    assign s_2_13_6 = s_12_13_7;
    assign s_1_13_6 = s_13_13_7;
    assign s_14_14_6 = s_1_14_7;
    assign s_13_14_6 = s_2_14_7;
    assign s_12_14_6 = s_3_14_7;
    assign s_11_14_6 = s_4_14_7;
    assign s_10_14_6 = s_5_14_7;
    assign s_9_14_6 = s_6_14_7;
    assign s_8_14_6 = s_7_14_7;
    assign s_7_14_6 = s_8_14_7;
    assign s_6_14_6 = s_9_14_7;
    assign s_5_14_6 = s_10_14_7;
    assign s_4_14_6 = s_11_14_7;
    assign s_3_14_6 = s_12_14_7;
    assign s_2_14_6 = s_13_14_7;
    assign s_1_14_6 = s_14_14_7;
    assign s_15_15_6 = s_1_15_7;
    assign s_14_15_6 = s_2_15_7;
    assign s_13_15_6 = s_3_15_7;
    assign s_12_15_6 = s_4_15_7;
    assign s_11_15_6 = s_5_15_7;
    assign s_10_15_6 = s_6_15_7;
    assign s_9_15_6 = s_7_15_7;
    assign s_8_15_6 = s_8_15_7;
    assign s_7_15_6 = s_9_15_7;
    assign s_6_15_6 = s_10_15_7;
    assign s_5_15_6 = s_11_15_7;
    assign s_4_15_6 = s_12_15_7;
    assign s_3_15_6 = s_13_15_7;
    assign s_2_15_6 = s_14_15_7;
    assign s_1_15_6 = s_15_15_7;
    assign s_16_16_6 = s_1_16_7;
    assign s_15_16_6 = s_2_16_7;
    assign s_14_16_6 = s_3_16_7;
    assign s_13_16_6 = s_4_16_7;
    assign s_12_16_6 = s_5_16_7;
    assign s_11_16_6 = s_6_16_7;
    assign s_10_16_6 = s_7_16_7;
    assign s_9_16_6 = s_8_16_7;
    assign s_8_16_6 = s_9_16_7;
    assign s_7_16_6 = s_10_16_7;
    assign s_6_16_6 = s_11_16_7;
    assign s_5_16_6 = s_12_16_7;
    assign s_4_16_6 = s_13_16_7;
    assign s_3_16_6 = s_14_16_7;
    assign s_2_16_6 = s_15_16_7;
    assign s_1_16_6 = s_16_16_7;
    assign s_17_17_6 = s_1_17_7;
    assign s_16_17_6 = s_2_17_7;
    assign s_15_17_6 = s_3_17_7;
    assign s_14_17_6 = s_4_17_7;
    assign s_13_17_6 = s_5_17_7;
    assign s_12_17_6 = s_6_17_7;
    assign s_11_17_6 = s_7_17_7;
    assign s_10_17_6 = s_8_17_7;
    assign s_9_17_6 = s_9_17_7;
    assign s_8_17_6 = s_10_17_7;
    assign s_7_17_6 = s_11_17_7;
    assign s_6_17_6 = s_12_17_7;
    assign s_5_17_6 = s_13_17_7;
    assign s_4_17_6 = s_14_17_7;
    assign s_3_17_6 = s_15_17_7;
    assign s_2_17_6 = s_16_17_7;
    assign s_1_17_6 = s_17_17_7;
    assign s_18_18_6 = s_1_18_7;
    assign s_17_18_6 = s_2_18_7;
    assign s_16_18_6 = s_3_18_7;
    assign s_15_18_6 = s_4_18_7;
    assign s_14_18_6 = s_5_18_7;
    assign s_13_18_6 = s_6_18_7;
    assign s_12_18_6 = s_7_18_7;
    assign s_11_18_6 = s_8_18_7;
    assign s_10_18_6 = s_9_18_7;
    assign s_9_18_6 = s_10_18_7;
    assign s_8_18_6 = s_11_18_7;
    assign s_7_18_6 = s_12_18_7;
    assign s_6_18_6 = s_13_18_7;
    assign s_5_18_6 = s_14_18_7;
    assign s_4_18_6 = s_15_18_7;
    assign s_3_18_6 = s_16_18_7;
    assign s_2_18_6 = s_17_18_7;
    assign s_1_18_6 = s_18_18_7;
    assign s_19_19_6 = s_1_19_7;
    assign s_18_19_6 = s_2_19_7;
    assign s_17_19_6 = s_3_19_7;
    assign s_16_19_6 = s_4_19_7;
    assign s_15_19_6 = s_5_19_7;
    assign s_14_19_6 = s_6_19_7;
    assign s_13_19_6 = s_7_19_7;
    assign s_12_19_6 = s_8_19_7;
    assign s_11_19_6 = s_9_19_7;
    assign s_10_19_6 = s_10_19_7;
    assign s_9_19_6 = s_11_19_7;
    assign s_8_19_6 = s_12_19_7;
    assign s_7_19_6 = s_13_19_7;
    assign s_6_19_6 = s_14_19_7;
    assign s_5_19_6 = s_15_19_7;
    assign s_4_19_6 = s_16_19_7;
    assign s_3_19_6 = s_17_19_7;
    assign s_2_19_6 = s_18_19_7;
    assign s_1_19_6 = s_19_19_7;
    HA HA4 (.A(s_1_20_7), .B(s_2_20_7), .S(s_19_20_6), .C(s_19_21_6));
    assign s_18_20_6 = s_3_20_7;
    assign s_17_20_6 = s_4_20_7;
    assign s_16_20_6 = s_5_20_7;
    assign s_15_20_6 = s_6_20_7;
    assign s_14_20_6 = s_7_20_7;
    assign s_13_20_6 = s_8_20_7;
    assign s_12_20_6 = s_9_20_7;
    assign s_11_20_6 = s_10_20_7;
    assign s_10_20_6 = s_11_20_7;
    assign s_9_20_6 = s_12_20_7;
    assign s_8_20_6 = s_13_20_7;
    assign s_7_20_6 = s_14_20_7;
    assign s_6_20_6 = s_15_20_7;
    assign s_5_20_6 = s_16_20_7;
    assign s_4_20_6 = s_17_20_7;
    assign s_3_20_6 = s_18_20_7;
    assign s_2_20_6 = s_19_20_7;
    assign s_1_20_6 = s_20_20_7;
    FA FA6 (.A(s_1_21_7), .B(s_2_21_7), .Cin(s_3_21_7), .S(s_18_21_6), .Cout(s_19_22_6));
    HA HA5 (.A(s_4_21_7), .B(s_5_21_7), .S(s_17_21_6), .C(s_18_22_6));
    assign s_16_21_6 = s_6_21_7;
    assign s_15_21_6 = s_7_21_7;
    assign s_14_21_6 = s_8_21_7;
    assign s_13_21_6 = s_9_21_7;
    assign s_12_21_6 = s_10_21_7;
    assign s_11_21_6 = s_11_21_7;
    assign s_10_21_6 = s_12_21_7;
    assign s_9_21_6 = s_13_21_7;
    assign s_8_21_6 = s_14_21_7;
    assign s_7_21_6 = s_15_21_7;
    assign s_6_21_6 = s_16_21_7;
    assign s_5_21_6 = s_17_21_7;
    assign s_4_21_6 = s_18_21_7;
    assign s_3_21_6 = s_19_21_7;
    assign s_2_21_6 = s_20_21_7;
    assign s_1_21_6 = s_21_21_7;
    FA FA7 (.A(s_1_22_7), .B(s_2_22_7), .Cin(s_3_22_7), .S(s_17_22_6), .Cout(s_19_23_6));
    FA FA8 (.A(s_4_22_7), .B(s_5_22_7), .Cin(s_6_22_7), .S(s_16_22_6), .Cout(s_18_23_6));
    HA HA6 (.A(s_7_22_7), .B(s_8_22_7), .S(s_15_22_6), .C(s_17_23_6));
    assign s_14_22_6 = s_9_22_7;
    assign s_13_22_6 = s_10_22_7;
    assign s_12_22_6 = s_11_22_7;
    assign s_11_22_6 = s_12_22_7;
    assign s_10_22_6 = s_13_22_7;
    assign s_9_22_6 = s_14_22_7;
    assign s_8_22_6 = s_15_22_7;
    assign s_7_22_6 = s_16_22_7;
    assign s_6_22_6 = s_17_22_7;
    assign s_5_22_6 = s_18_22_7;
    assign s_4_22_6 = s_19_22_7;
    assign s_3_22_6 = s_20_22_7;
    assign s_2_22_6 = s_21_22_7;
    assign s_1_22_6 = s_22_22_7;
    FA FA9 (.A(s_1_23_7), .B(s_2_23_7), .Cin(s_3_23_7), .S(s_16_23_6), .Cout(s_19_24_6));
    FA FA10 (.A(s_4_23_7), .B(s_5_23_7), .Cin(s_6_23_7), .S(s_15_23_6), .Cout(s_18_24_6));
    FA FA11 (.A(s_7_23_7), .B(s_8_23_7), .Cin(s_9_23_7), .S(s_14_23_6), .Cout(s_17_24_6));
    HA HA7 (.A(s_10_23_7), .B(s_11_23_7), .S(s_13_23_6), .C(s_16_24_6));
    assign s_12_23_6 = s_12_23_7;
    assign s_11_23_6 = s_13_23_7;
    assign s_10_23_6 = s_14_23_7;
    assign s_9_23_6 = s_15_23_7;
    assign s_8_23_6 = s_16_23_7;
    assign s_7_23_6 = s_17_23_7;
    assign s_6_23_6 = s_18_23_7;
    assign s_5_23_6 = s_19_23_7;
    assign s_4_23_6 = s_20_23_7;
    assign s_3_23_6 = s_21_23_7;
    assign s_2_23_6 = s_22_23_7;
    assign s_1_23_6 = s_23_23_7;
    FA FA12 (.A(s_1_24_7), .B(s_2_24_7), .Cin(s_3_24_7), .S(s_15_24_6), .Cout(s_19_25_6));
    FA FA13 (.A(s_4_24_7), .B(s_5_24_7), .Cin(s_6_24_7), .S(s_14_24_6), .Cout(s_18_25_6));
    FA FA14 (.A(s_7_24_7), .B(s_8_24_7), .Cin(s_9_24_7), .S(s_13_24_6), .Cout(s_17_25_6));
    FA FA15 (.A(s_10_24_7), .B(s_11_24_7), .Cin(s_12_24_7), .S(s_12_24_6), .Cout(s_16_25_6));
    HA HA8 (.A(s_13_24_7), .B(s_14_24_7), .S(s_11_24_6), .C(s_15_25_6));
    assign s_10_24_6 = s_15_24_7;
    assign s_9_24_6 = s_16_24_7;
    assign s_8_24_6 = s_17_24_7;
    assign s_7_24_6 = s_18_24_7;
    assign s_6_24_6 = s_19_24_7;
    assign s_5_24_6 = s_20_24_7;
    assign s_4_24_6 = s_21_24_7;
    assign s_3_24_6 = s_22_24_7;
    assign s_2_24_6 = s_23_24_7;
    assign s_1_24_6 = s_24_24_7;
    FA FA16 (.A(s_1_25_7), .B(s_2_25_7), .Cin(s_3_25_7), .S(s_14_25_6), .Cout(s_19_26_6));
    FA FA17 (.A(s_4_25_7), .B(s_5_25_7), .Cin(s_6_25_7), .S(s_13_25_6), .Cout(s_18_26_6));
    FA FA18 (.A(s_7_25_7), .B(s_8_25_7), .Cin(s_9_25_7), .S(s_12_25_6), .Cout(s_17_26_6));
    FA FA19 (.A(s_10_25_7), .B(s_11_25_7), .Cin(s_12_25_7), .S(s_11_25_6), .Cout(s_16_26_6));
    FA FA20 (.A(s_13_25_7), .B(s_14_25_7), .Cin(s_15_25_7), .S(s_10_25_6), .Cout(s_15_26_6));
    HA HA9 (.A(s_16_25_7), .B(s_17_25_7), .S(s_9_25_6), .C(s_14_26_6));
    assign s_8_25_6 = s_18_25_7;
    assign s_7_25_6 = s_19_25_7;
    assign s_6_25_6 = s_20_25_7;
    assign s_5_25_6 = s_21_25_7;
    assign s_4_25_6 = s_22_25_7;
    assign s_3_25_6 = s_23_25_7;
    assign s_2_25_6 = s_24_25_7;
    assign s_1_25_6 = s_25_25_7;
    FA FA21 (.A(s_1_26_7), .B(s_2_26_7), .Cin(s_3_26_7), .S(s_13_26_6), .Cout(s_19_27_6));
    FA FA22 (.A(s_4_26_7), .B(s_5_26_7), .Cin(s_6_26_7), .S(s_12_26_6), .Cout(s_18_27_6));
    FA FA23 (.A(s_7_26_7), .B(s_8_26_7), .Cin(s_9_26_7), .S(s_11_26_6), .Cout(s_17_27_6));
    FA FA24 (.A(s_10_26_7), .B(s_11_26_7), .Cin(s_12_26_7), .S(s_10_26_6), .Cout(s_16_27_6));
    FA FA25 (.A(s_13_26_7), .B(s_14_26_7), .Cin(s_15_26_7), .S(s_9_26_6), .Cout(s_15_27_6));
    FA FA26 (.A(s_16_26_7), .B(s_17_26_7), .Cin(s_18_26_7), .S(s_8_26_6), .Cout(s_14_27_6));
    HA HA10 (.A(s_19_26_7), .B(s_20_26_7), .S(s_7_26_6), .C(s_13_27_6));
    assign s_6_26_6 = s_21_26_7;
    assign s_5_26_6 = s_22_26_7;
    assign s_4_26_6 = s_23_26_7;
    assign s_3_26_6 = s_24_26_7;
    assign s_2_26_6 = s_25_26_7;
    assign s_1_26_6 = s_26_26_7;
    FA FA27 (.A(s_1_27_7), .B(s_2_27_7), .Cin(s_3_27_7), .S(s_12_27_6), .Cout(s_19_28_6));
    FA FA28 (.A(s_4_27_7), .B(s_5_27_7), .Cin(s_6_27_7), .S(s_11_27_6), .Cout(s_18_28_6));
    FA FA29 (.A(s_7_27_7), .B(s_8_27_7), .Cin(s_9_27_7), .S(s_10_27_6), .Cout(s_17_28_6));
    FA FA30 (.A(s_10_27_7), .B(s_11_27_7), .Cin(s_12_27_7), .S(s_9_27_6), .Cout(s_16_28_6));
    FA FA31 (.A(s_13_27_7), .B(s_14_27_7), .Cin(s_15_27_7), .S(s_8_27_6), .Cout(s_15_28_6));
    FA FA32 (.A(s_16_27_7), .B(s_17_27_7), .Cin(s_18_27_7), .S(s_7_27_6), .Cout(s_14_28_6));
    FA FA33 (.A(s_19_27_7), .B(s_20_27_7), .Cin(s_21_27_7), .S(s_6_27_6), .Cout(s_13_28_6));
    HA HA11 (.A(s_22_27_7), .B(s_23_27_7), .S(s_5_27_6), .C(s_12_28_6));
    assign s_4_27_6 = s_24_27_7;
    assign s_3_27_6 = s_25_27_7;
    assign s_2_27_6 = s_26_27_7;
    assign s_1_27_6 = s_27_27_7;
    FA FA34 (.A(s_1_28_7), .B(s_2_28_7), .Cin(s_3_28_7), .S(s_11_28_6), .Cout(s_19_29_6));
    FA FA35 (.A(s_4_28_7), .B(s_5_28_7), .Cin(s_6_28_7), .S(s_10_28_6), .Cout(s_18_29_6));
    FA FA36 (.A(s_7_28_7), .B(s_8_28_7), .Cin(s_9_28_7), .S(s_9_28_6), .Cout(s_17_29_6));
    FA FA37 (.A(s_10_28_7), .B(s_11_28_7), .Cin(s_12_28_7), .S(s_8_28_6), .Cout(s_16_29_6));
    FA FA38 (.A(s_13_28_7), .B(s_14_28_7), .Cin(s_15_28_7), .S(s_7_28_6), .Cout(s_15_29_6));
    FA FA39 (.A(s_16_28_7), .B(s_17_28_7), .Cin(s_18_28_7), .S(s_6_28_6), .Cout(s_14_29_6));
    FA FA40 (.A(s_19_28_7), .B(s_20_28_7), .Cin(s_21_28_7), .S(s_5_28_6), .Cout(s_13_29_6));
    FA FA41 (.A(s_22_28_7), .B(s_23_28_7), .Cin(s_24_28_7), .S(s_4_28_6), .Cout(s_12_29_6));
    HA HA12 (.A(s_25_28_7), .B(s_26_28_7), .S(s_3_28_6), .C(s_11_29_6));
    assign s_2_28_6 = s_27_28_7;
    assign s_1_28_6 = s_28_28_7;
    FA FA42 (.A(s_1_29_7), .B(s_2_29_7), .Cin(s_3_29_7), .S(s_10_29_6), .Cout(s_19_30_6));
    FA FA43 (.A(s_4_29_7), .B(s_5_29_7), .Cin(s_6_29_7), .S(s_9_29_6), .Cout(s_18_30_6));
    FA FA44 (.A(s_7_29_7), .B(s_8_29_7), .Cin(s_9_29_7), .S(s_8_29_6), .Cout(s_17_30_6));
    FA FA45 (.A(s_10_29_7), .B(s_11_29_7), .Cin(s_12_29_7), .S(s_7_29_6), .Cout(s_16_30_6));
    FA FA46 (.A(s_13_29_7), .B(s_14_29_7), .Cin(s_15_29_7), .S(s_6_29_6), .Cout(s_15_30_6));
    FA FA47 (.A(s_16_29_7), .B(s_17_29_7), .Cin(s_18_29_7), .S(s_5_29_6), .Cout(s_14_30_6));
    FA FA48 (.A(s_19_29_7), .B(s_20_29_7), .Cin(s_21_29_7), .S(s_4_29_6), .Cout(s_13_30_6));
    FA FA49 (.A(s_22_29_7), .B(s_23_29_7), .Cin(s_24_29_7), .S(s_3_29_6), .Cout(s_12_30_6));
    FA FA50 (.A(s_25_29_7), .B(s_26_29_7), .Cin(s_27_29_7), .S(s_2_29_6), .Cout(s_11_30_6));
    assign s_1_29_6 = s_28_29_7;
    FA FA51 (.A(s_1_30_7), .B(s_2_30_7), .Cin(s_3_30_7), .S(s_10_30_6), .Cout(s_19_31_6));
    FA FA52 (.A(s_4_30_7), .B(s_5_30_7), .Cin(s_6_30_7), .S(s_9_30_6), .Cout(s_18_31_6));
    FA FA53 (.A(s_7_30_7), .B(s_8_30_7), .Cin(s_9_30_7), .S(s_8_30_6), .Cout(s_17_31_6));
    FA FA54 (.A(s_10_30_7), .B(s_11_30_7), .Cin(s_12_30_7), .S(s_7_30_6), .Cout(s_16_31_6));
    FA FA55 (.A(s_13_30_7), .B(s_14_30_7), .Cin(s_15_30_7), .S(s_6_30_6), .Cout(s_15_31_6));
    FA FA56 (.A(s_16_30_7), .B(s_17_30_7), .Cin(s_18_30_7), .S(s_5_30_6), .Cout(s_14_31_6));
    FA FA57 (.A(s_19_30_7), .B(s_20_30_7), .Cin(s_21_30_7), .S(s_4_30_6), .Cout(s_13_31_6));
    FA FA58 (.A(s_22_30_7), .B(s_23_30_7), .Cin(s_24_30_7), .S(s_3_30_6), .Cout(s_12_31_6));
    FA FA59 (.A(s_25_30_7), .B(s_26_30_7), .Cin(s_27_30_7), .S(s_2_30_6), .Cout(s_11_31_6));
    assign s_1_30_6 = s_28_30_7;
    FA FA60 (.A(s_1_31_7), .B(s_2_31_7), .Cin(s_3_31_7), .S(s_10_31_6), .Cout(s_19_32_6));
    FA FA61 (.A(s_4_31_7), .B(s_5_31_7), .Cin(s_6_31_7), .S(s_9_31_6), .Cout(s_18_32_6));
    FA FA62 (.A(s_7_31_7), .B(s_8_31_7), .Cin(s_9_31_7), .S(s_8_31_6), .Cout(s_17_32_6));
    FA FA63 (.A(s_10_31_7), .B(s_11_31_7), .Cin(s_12_31_7), .S(s_7_31_6), .Cout(s_16_32_6));
    FA FA64 (.A(s_13_31_7), .B(s_14_31_7), .Cin(s_15_31_7), .S(s_6_31_6), .Cout(s_15_32_6));
    FA FA65 (.A(s_16_31_7), .B(s_17_31_7), .Cin(s_18_31_7), .S(s_5_31_6), .Cout(s_14_32_6));
    FA FA66 (.A(s_19_31_7), .B(s_20_31_7), .Cin(s_21_31_7), .S(s_4_31_6), .Cout(s_13_32_6));
    FA FA67 (.A(s_22_31_7), .B(s_23_31_7), .Cin(s_24_31_7), .S(s_3_31_6), .Cout(s_12_32_6));
    FA FA68 (.A(s_25_31_7), .B(s_26_31_7), .Cin(s_27_31_7), .S(s_2_31_6), .Cout(s_11_32_6));
    assign s_1_31_6 = s_28_31_7;
    FA FA69 (.A(s_1_32_7), .B(s_2_32_7), .Cin(s_3_32_7), .S(s_10_32_6), .Cout(s_19_33_6));
    FA FA70 (.A(s_4_32_7), .B(s_5_32_7), .Cin(s_6_32_7), .S(s_9_32_6), .Cout(s_18_33_6));
    FA FA71 (.A(s_7_32_7), .B(s_8_32_7), .Cin(s_9_32_7), .S(s_8_32_6), .Cout(s_17_33_6));
    FA FA72 (.A(s_10_32_7), .B(s_11_32_7), .Cin(s_12_32_7), .S(s_7_32_6), .Cout(s_16_33_6));
    FA FA73 (.A(s_13_32_7), .B(s_14_32_7), .Cin(s_15_32_7), .S(s_6_32_6), .Cout(s_15_33_6));
    FA FA74 (.A(s_16_32_7), .B(s_17_32_7), .Cin(s_18_32_7), .S(s_5_32_6), .Cout(s_14_33_6));
    FA FA75 (.A(s_19_32_7), .B(s_20_32_7), .Cin(s_21_32_7), .S(s_4_32_6), .Cout(s_13_33_6));
    FA FA76 (.A(s_22_32_7), .B(s_23_32_7), .Cin(s_24_32_7), .S(s_3_32_6), .Cout(s_12_33_6));
    FA FA77 (.A(s_25_32_7), .B(s_26_32_7), .Cin(s_27_32_7), .S(s_2_32_6), .Cout(s_11_33_6));
    assign s_1_32_6 = s_28_32_7;
    // total 9 half adders and 72 full adders
    // d_7 = 19 done

    assign s_1_1_5 = s_1_1_6;
    assign s_2_2_5 = s_1_2_6;
    assign s_1_2_5 = s_2_2_6;
    assign s_3_3_5 = s_1_3_6;
    assign s_2_3_5 = s_2_3_6;
    assign s_1_3_5 = s_3_3_6;
    assign s_4_4_5 = s_1_4_6;
    assign s_3_4_5 = s_2_4_6;
    assign s_2_4_5 = s_3_4_6;
    assign s_1_4_5 = s_4_4_6;
    assign s_5_5_5 = s_1_5_6;
    assign s_4_5_5 = s_2_5_6;
    assign s_3_5_5 = s_3_5_6;
    assign s_2_5_5 = s_4_5_6;
    assign s_1_5_5 = s_5_5_6;
    assign s_6_6_5 = s_1_6_6;
    assign s_5_6_5 = s_2_6_6;
    assign s_4_6_5 = s_3_6_6;
    assign s_3_6_5 = s_4_6_6;
    assign s_2_6_5 = s_5_6_6;
    assign s_1_6_5 = s_6_6_6;
    assign s_7_7_5 = s_1_7_6;
    assign s_6_7_5 = s_2_7_6;
    assign s_5_7_5 = s_3_7_6;
    assign s_4_7_5 = s_4_7_6;
    assign s_3_7_5 = s_5_7_6;
    assign s_2_7_5 = s_6_7_6;
    assign s_1_7_5 = s_7_7_6;
    assign s_8_8_5 = s_1_8_6;
    assign s_7_8_5 = s_2_8_6;
    assign s_6_8_5 = s_3_8_6;
    assign s_5_8_5 = s_4_8_6;
    assign s_4_8_5 = s_5_8_6;
    assign s_3_8_5 = s_6_8_6;
    assign s_2_8_5 = s_7_8_6;
    assign s_1_8_5 = s_8_8_6;
    assign s_9_9_5 = s_1_9_6;
    assign s_8_9_5 = s_2_9_6;
    assign s_7_9_5 = s_3_9_6;
    assign s_6_9_5 = s_4_9_6;
    assign s_5_9_5 = s_5_9_6;
    assign s_4_9_5 = s_6_9_6;
    assign s_3_9_5 = s_7_9_6;
    assign s_2_9_5 = s_8_9_6;
    assign s_1_9_5 = s_9_9_6;
    assign s_10_10_5 = s_1_10_6;
    assign s_9_10_5 = s_2_10_6;
    assign s_8_10_5 = s_3_10_6;
    assign s_7_10_5 = s_4_10_6;
    assign s_6_10_5 = s_5_10_6;
    assign s_5_10_5 = s_6_10_6;
    assign s_4_10_5 = s_7_10_6;
    assign s_3_10_5 = s_8_10_6;
    assign s_2_10_5 = s_9_10_6;
    assign s_1_10_5 = s_10_10_6;
    assign s_11_11_5 = s_1_11_6;
    assign s_10_11_5 = s_2_11_6;
    assign s_9_11_5 = s_3_11_6;
    assign s_8_11_5 = s_4_11_6;
    assign s_7_11_5 = s_5_11_6;
    assign s_6_11_5 = s_6_11_6;
    assign s_5_11_5 = s_7_11_6;
    assign s_4_11_5 = s_8_11_6;
    assign s_3_11_5 = s_9_11_6;
    assign s_2_11_5 = s_10_11_6;
    assign s_1_11_5 = s_11_11_6;
    assign s_12_12_5 = s_1_12_6;
    assign s_11_12_5 = s_2_12_6;
    assign s_10_12_5 = s_3_12_6;
    assign s_9_12_5 = s_4_12_6;
    assign s_8_12_5 = s_5_12_6;
    assign s_7_12_5 = s_6_12_6;
    assign s_6_12_5 = s_7_12_6;
    assign s_5_12_5 = s_8_12_6;
    assign s_4_12_5 = s_9_12_6;
    assign s_3_12_5 = s_10_12_6;
    assign s_2_12_5 = s_11_12_6;
    assign s_1_12_5 = s_12_12_6;
    assign s_13_13_5 = s_1_13_6;
    assign s_12_13_5 = s_2_13_6;
    assign s_11_13_5 = s_3_13_6;
    assign s_10_13_5 = s_4_13_6;
    assign s_9_13_5 = s_5_13_6;
    assign s_8_13_5 = s_6_13_6;
    assign s_7_13_5 = s_7_13_6;
    assign s_6_13_5 = s_8_13_6;
    assign s_5_13_5 = s_9_13_6;
    assign s_4_13_5 = s_10_13_6;
    assign s_3_13_5 = s_11_13_6;
    assign s_2_13_5 = s_12_13_6;
    assign s_1_13_5 = s_13_13_6;
    HA HA13 (.A(s_1_14_6), .B(s_2_14_6), .S(s_13_14_5), .C(s_13_15_5));
    assign s_12_14_5 = s_3_14_6;
    assign s_11_14_5 = s_4_14_6;
    assign s_10_14_5 = s_5_14_6;
    assign s_9_14_5 = s_6_14_6;
    assign s_8_14_5 = s_7_14_6;
    assign s_7_14_5 = s_8_14_6;
    assign s_6_14_5 = s_9_14_6;
    assign s_5_14_5 = s_10_14_6;
    assign s_4_14_5 = s_11_14_6;
    assign s_3_14_5 = s_12_14_6;
    assign s_2_14_5 = s_13_14_6;
    assign s_1_14_5 = s_14_14_6;
    FA FA78 (.A(s_1_15_6), .B(s_2_15_6), .Cin(s_3_15_6), .S(s_12_15_5), .Cout(s_13_16_5));
    HA HA14 (.A(s_4_15_6), .B(s_5_15_6), .S(s_11_15_5), .C(s_12_16_5));
    assign s_10_15_5 = s_6_15_6;
    assign s_9_15_5 = s_7_15_6;
    assign s_8_15_5 = s_8_15_6;
    assign s_7_15_5 = s_9_15_6;
    assign s_6_15_5 = s_10_15_6;
    assign s_5_15_5 = s_11_15_6;
    assign s_4_15_5 = s_12_15_6;
    assign s_3_15_5 = s_13_15_6;
    assign s_2_15_5 = s_14_15_6;
    assign s_1_15_5 = s_15_15_6;
    FA FA79 (.A(s_1_16_6), .B(s_2_16_6), .Cin(s_3_16_6), .S(s_11_16_5), .Cout(s_13_17_5));
    FA FA80 (.A(s_4_16_6), .B(s_5_16_6), .Cin(s_6_16_6), .S(s_10_16_5), .Cout(s_12_17_5));
    HA HA15 (.A(s_7_16_6), .B(s_8_16_6), .S(s_9_16_5), .C(s_11_17_5));
    assign s_8_16_5 = s_9_16_6;
    assign s_7_16_5 = s_10_16_6;
    assign s_6_16_5 = s_11_16_6;
    assign s_5_16_5 = s_12_16_6;
    assign s_4_16_5 = s_13_16_6;
    assign s_3_16_5 = s_14_16_6;
    assign s_2_16_5 = s_15_16_6;
    assign s_1_16_5 = s_16_16_6;
    FA FA81 (.A(s_1_17_6), .B(s_2_17_6), .Cin(s_3_17_6), .S(s_10_17_5), .Cout(s_13_18_5));
    FA FA82 (.A(s_4_17_6), .B(s_5_17_6), .Cin(s_6_17_6), .S(s_9_17_5), .Cout(s_12_18_5));
    FA FA83 (.A(s_7_17_6), .B(s_8_17_6), .Cin(s_9_17_6), .S(s_8_17_5), .Cout(s_11_18_5));
    HA HA16 (.A(s_10_17_6), .B(s_11_17_6), .S(s_7_17_5), .C(s_10_18_5));
    assign s_6_17_5 = s_12_17_6;
    assign s_5_17_5 = s_13_17_6;
    assign s_4_17_5 = s_14_17_6;
    assign s_3_17_5 = s_15_17_6;
    assign s_2_17_5 = s_16_17_6;
    assign s_1_17_5 = s_17_17_6;
    FA FA84 (.A(s_1_18_6), .B(s_2_18_6), .Cin(s_3_18_6), .S(s_9_18_5), .Cout(s_13_19_5));
    FA FA85 (.A(s_4_18_6), .B(s_5_18_6), .Cin(s_6_18_6), .S(s_8_18_5), .Cout(s_12_19_5));
    FA FA86 (.A(s_7_18_6), .B(s_8_18_6), .Cin(s_9_18_6), .S(s_7_18_5), .Cout(s_11_19_5));
    FA FA87 (.A(s_10_18_6), .B(s_11_18_6), .Cin(s_12_18_6), .S(s_6_18_5), .Cout(s_10_19_5));
    HA HA17 (.A(s_13_18_6), .B(s_14_18_6), .S(s_5_18_5), .C(s_9_19_5));
    assign s_4_18_5 = s_15_18_6;
    assign s_3_18_5 = s_16_18_6;
    assign s_2_18_5 = s_17_18_6;
    assign s_1_18_5 = s_18_18_6;
    FA FA88 (.A(s_1_19_6), .B(s_2_19_6), .Cin(s_3_19_6), .S(s_8_19_5), .Cout(s_13_20_5));
    FA FA89 (.A(s_4_19_6), .B(s_5_19_6), .Cin(s_6_19_6), .S(s_7_19_5), .Cout(s_12_20_5));
    FA FA90 (.A(s_7_19_6), .B(s_8_19_6), .Cin(s_9_19_6), .S(s_6_19_5), .Cout(s_11_20_5));
    FA FA91 (.A(s_10_19_6), .B(s_11_19_6), .Cin(s_12_19_6), .S(s_5_19_5), .Cout(s_10_20_5));
    FA FA92 (.A(s_13_19_6), .B(s_14_19_6), .Cin(s_15_19_6), .S(s_4_19_5), .Cout(s_9_20_5));
    HA HA18 (.A(s_16_19_6), .B(s_17_19_6), .S(s_3_19_5), .C(s_8_20_5));
    assign s_2_19_5 = s_18_19_6;
    assign s_1_19_5 = s_19_19_6;
    FA FA93 (.A(s_1_20_6), .B(s_2_20_6), .Cin(s_3_20_6), .S(s_7_20_5), .Cout(s_13_21_5));
    FA FA94 (.A(s_4_20_6), .B(s_5_20_6), .Cin(s_6_20_6), .S(s_6_20_5), .Cout(s_12_21_5));
    FA FA95 (.A(s_7_20_6), .B(s_8_20_6), .Cin(s_9_20_6), .S(s_5_20_5), .Cout(s_11_21_5));
    FA FA96 (.A(s_10_20_6), .B(s_11_20_6), .Cin(s_12_20_6), .S(s_4_20_5), .Cout(s_10_21_5));
    FA FA97 (.A(s_13_20_6), .B(s_14_20_6), .Cin(s_15_20_6), .S(s_3_20_5), .Cout(s_9_21_5));
    FA FA98 (.A(s_16_20_6), .B(s_17_20_6), .Cin(s_18_20_6), .S(s_2_20_5), .Cout(s_8_21_5));
    assign s_1_20_5 = s_19_20_6;
    FA FA99 (.A(s_1_21_6), .B(s_2_21_6), .Cin(s_3_21_6), .S(s_7_21_5), .Cout(s_13_22_5));
    FA FA100 (.A(s_4_21_6), .B(s_5_21_6), .Cin(s_6_21_6), .S(s_6_21_5), .Cout(s_12_22_5));
    FA FA101 (.A(s_7_21_6), .B(s_8_21_6), .Cin(s_9_21_6), .S(s_5_21_5), .Cout(s_11_22_5));
    FA FA102 (.A(s_10_21_6), .B(s_11_21_6), .Cin(s_12_21_6), .S(s_4_21_5), .Cout(s_10_22_5));
    FA FA103 (.A(s_13_21_6), .B(s_14_21_6), .Cin(s_15_21_6), .S(s_3_21_5), .Cout(s_9_22_5));
    FA FA104 (.A(s_16_21_6), .B(s_17_21_6), .Cin(s_18_21_6), .S(s_2_21_5), .Cout(s_8_22_5));
    assign s_1_21_5 = s_19_21_6;
    FA FA105 (.A(s_1_22_6), .B(s_2_22_6), .Cin(s_3_22_6), .S(s_7_22_5), .Cout(s_13_23_5));
    FA FA106 (.A(s_4_22_6), .B(s_5_22_6), .Cin(s_6_22_6), .S(s_6_22_5), .Cout(s_12_23_5));
    FA FA107 (.A(s_7_22_6), .B(s_8_22_6), .Cin(s_9_22_6), .S(s_5_22_5), .Cout(s_11_23_5));
    FA FA108 (.A(s_10_22_6), .B(s_11_22_6), .Cin(s_12_22_6), .S(s_4_22_5), .Cout(s_10_23_5));
    FA FA109 (.A(s_13_22_6), .B(s_14_22_6), .Cin(s_15_22_6), .S(s_3_22_5), .Cout(s_9_23_5));
    FA FA110 (.A(s_16_22_6), .B(s_17_22_6), .Cin(s_18_22_6), .S(s_2_22_5), .Cout(s_8_23_5));
    assign s_1_22_5 = s_19_22_6;
    FA FA111 (.A(s_1_23_6), .B(s_2_23_6), .Cin(s_3_23_6), .S(s_7_23_5), .Cout(s_13_24_5));
    FA FA112 (.A(s_4_23_6), .B(s_5_23_6), .Cin(s_6_23_6), .S(s_6_23_5), .Cout(s_12_24_5));
    FA FA113 (.A(s_7_23_6), .B(s_8_23_6), .Cin(s_9_23_6), .S(s_5_23_5), .Cout(s_11_24_5));
    FA FA114 (.A(s_10_23_6), .B(s_11_23_6), .Cin(s_12_23_6), .S(s_4_23_5), .Cout(s_10_24_5));
    FA FA115 (.A(s_13_23_6), .B(s_14_23_6), .Cin(s_15_23_6), .S(s_3_23_5), .Cout(s_9_24_5));
    FA FA116 (.A(s_16_23_6), .B(s_17_23_6), .Cin(s_18_23_6), .S(s_2_23_5), .Cout(s_8_24_5));
    assign s_1_23_5 = s_19_23_6;
    FA FA117 (.A(s_1_24_6), .B(s_2_24_6), .Cin(s_3_24_6), .S(s_7_24_5), .Cout(s_13_25_5));
    FA FA118 (.A(s_4_24_6), .B(s_5_24_6), .Cin(s_6_24_6), .S(s_6_24_5), .Cout(s_12_25_5));
    FA FA119 (.A(s_7_24_6), .B(s_8_24_6), .Cin(s_9_24_6), .S(s_5_24_5), .Cout(s_11_25_5));
    FA FA120 (.A(s_10_24_6), .B(s_11_24_6), .Cin(s_12_24_6), .S(s_4_24_5), .Cout(s_10_25_5));
    FA FA121 (.A(s_13_24_6), .B(s_14_24_6), .Cin(s_15_24_6), .S(s_3_24_5), .Cout(s_9_25_5));
    FA FA122 (.A(s_16_24_6), .B(s_17_24_6), .Cin(s_18_24_6), .S(s_2_24_5), .Cout(s_8_25_5));
    assign s_1_24_5 = s_19_24_6;
    FA FA123 (.A(s_1_25_6), .B(s_2_25_6), .Cin(s_3_25_6), .S(s_7_25_5), .Cout(s_13_26_5));
    FA FA124 (.A(s_4_25_6), .B(s_5_25_6), .Cin(s_6_25_6), .S(s_6_25_5), .Cout(s_12_26_5));
    FA FA125 (.A(s_7_25_6), .B(s_8_25_6), .Cin(s_9_25_6), .S(s_5_25_5), .Cout(s_11_26_5));
    FA FA126 (.A(s_10_25_6), .B(s_11_25_6), .Cin(s_12_25_6), .S(s_4_25_5), .Cout(s_10_26_5));
    FA FA127 (.A(s_13_25_6), .B(s_14_25_6), .Cin(s_15_25_6), .S(s_3_25_5), .Cout(s_9_26_5));
    FA FA128 (.A(s_16_25_6), .B(s_17_25_6), .Cin(s_18_25_6), .S(s_2_25_5), .Cout(s_8_26_5));
    assign s_1_25_5 = s_19_25_6;
    FA FA129 (.A(s_1_26_6), .B(s_2_26_6), .Cin(s_3_26_6), .S(s_7_26_5), .Cout(s_13_27_5));
    FA FA130 (.A(s_4_26_6), .B(s_5_26_6), .Cin(s_6_26_6), .S(s_6_26_5), .Cout(s_12_27_5));
    FA FA131 (.A(s_7_26_6), .B(s_8_26_6), .Cin(s_9_26_6), .S(s_5_26_5), .Cout(s_11_27_5));
    FA FA132 (.A(s_10_26_6), .B(s_11_26_6), .Cin(s_12_26_6), .S(s_4_26_5), .Cout(s_10_27_5));
    FA FA133 (.A(s_13_26_6), .B(s_14_26_6), .Cin(s_15_26_6), .S(s_3_26_5), .Cout(s_9_27_5));
    FA FA134 (.A(s_16_26_6), .B(s_17_26_6), .Cin(s_18_26_6), .S(s_2_26_5), .Cout(s_8_27_5));
    assign s_1_26_5 = s_19_26_6;
    FA FA135 (.A(s_1_27_6), .B(s_2_27_6), .Cin(s_3_27_6), .S(s_7_27_5), .Cout(s_13_28_5));
    FA FA136 (.A(s_4_27_6), .B(s_5_27_6), .Cin(s_6_27_6), .S(s_6_27_5), .Cout(s_12_28_5));
    FA FA137 (.A(s_7_27_6), .B(s_8_27_6), .Cin(s_9_27_6), .S(s_5_27_5), .Cout(s_11_28_5));
    FA FA138 (.A(s_10_27_6), .B(s_11_27_6), .Cin(s_12_27_6), .S(s_4_27_5), .Cout(s_10_28_5));
    FA FA139 (.A(s_13_27_6), .B(s_14_27_6), .Cin(s_15_27_6), .S(s_3_27_5), .Cout(s_9_28_5));
    FA FA140 (.A(s_16_27_6), .B(s_17_27_6), .Cin(s_18_27_6), .S(s_2_27_5), .Cout(s_8_28_5));
    assign s_1_27_5 = s_19_27_6;
    FA FA141 (.A(s_1_28_6), .B(s_2_28_6), .Cin(s_3_28_6), .S(s_7_28_5), .Cout(s_13_29_5));
    FA FA142 (.A(s_4_28_6), .B(s_5_28_6), .Cin(s_6_28_6), .S(s_6_28_5), .Cout(s_12_29_5));
    FA FA143 (.A(s_7_28_6), .B(s_8_28_6), .Cin(s_9_28_6), .S(s_5_28_5), .Cout(s_11_29_5));
    FA FA144 (.A(s_10_28_6), .B(s_11_28_6), .Cin(s_12_28_6), .S(s_4_28_5), .Cout(s_10_29_5));
    FA FA145 (.A(s_13_28_6), .B(s_14_28_6), .Cin(s_15_28_6), .S(s_3_28_5), .Cout(s_9_29_5));
    FA FA146 (.A(s_16_28_6), .B(s_17_28_6), .Cin(s_18_28_6), .S(s_2_28_5), .Cout(s_8_29_5));
    assign s_1_28_5 = s_19_28_6;
    FA FA147 (.A(s_1_29_6), .B(s_2_29_6), .Cin(s_3_29_6), .S(s_7_29_5), .Cout(s_13_30_5));
    FA FA148 (.A(s_4_29_6), .B(s_5_29_6), .Cin(s_6_29_6), .S(s_6_29_5), .Cout(s_12_30_5));
    FA FA149 (.A(s_7_29_6), .B(s_8_29_6), .Cin(s_9_29_6), .S(s_5_29_5), .Cout(s_11_30_5));
    FA FA150 (.A(s_10_29_6), .B(s_11_29_6), .Cin(s_12_29_6), .S(s_4_29_5), .Cout(s_10_30_5));
    FA FA151 (.A(s_13_29_6), .B(s_14_29_6), .Cin(s_15_29_6), .S(s_3_29_5), .Cout(s_9_30_5));
    FA FA152 (.A(s_16_29_6), .B(s_17_29_6), .Cin(s_18_29_6), .S(s_2_29_5), .Cout(s_8_30_5));
    assign s_1_29_5 = s_19_29_6;
    FA FA153 (.A(s_1_30_6), .B(s_2_30_6), .Cin(s_3_30_6), .S(s_7_30_5), .Cout(s_13_31_5));
    FA FA154 (.A(s_4_30_6), .B(s_5_30_6), .Cin(s_6_30_6), .S(s_6_30_5), .Cout(s_12_31_5));
    FA FA155 (.A(s_7_30_6), .B(s_8_30_6), .Cin(s_9_30_6), .S(s_5_30_5), .Cout(s_11_31_5));
    FA FA156 (.A(s_10_30_6), .B(s_11_30_6), .Cin(s_12_30_6), .S(s_4_30_5), .Cout(s_10_31_5));
    FA FA157 (.A(s_13_30_6), .B(s_14_30_6), .Cin(s_15_30_6), .S(s_3_30_5), .Cout(s_9_31_5));
    FA FA158 (.A(s_16_30_6), .B(s_17_30_6), .Cin(s_18_30_6), .S(s_2_30_5), .Cout(s_8_31_5));
    assign s_1_30_5 = s_19_30_6;
    FA FA159 (.A(s_1_31_6), .B(s_2_31_6), .Cin(s_3_31_6), .S(s_7_31_5), .Cout(s_13_32_5));
    FA FA160 (.A(s_4_31_6), .B(s_5_31_6), .Cin(s_6_31_6), .S(s_6_31_5), .Cout(s_12_32_5));
    FA FA161 (.A(s_7_31_6), .B(s_8_31_6), .Cin(s_9_31_6), .S(s_5_31_5), .Cout(s_11_32_5));
    FA FA162 (.A(s_10_31_6), .B(s_11_31_6), .Cin(s_12_31_6), .S(s_4_31_5), .Cout(s_10_32_5));
    FA FA163 (.A(s_13_31_6), .B(s_14_31_6), .Cin(s_15_31_6), .S(s_3_31_5), .Cout(s_9_32_5));
    FA FA164 (.A(s_16_31_6), .B(s_17_31_6), .Cin(s_18_31_6), .S(s_2_31_5), .Cout(s_8_32_5));
    assign s_1_31_5 = s_19_31_6;
    FA FA165 (.A(s_1_32_6), .B(s_2_32_6), .Cin(s_3_32_6), .S(s_7_32_5), .Cout(s_13_33_5));
    FA FA166 (.A(s_4_32_6), .B(s_5_32_6), .Cin(s_6_32_6), .S(s_6_32_5), .Cout(s_12_33_5));
    FA FA167 (.A(s_7_32_6), .B(s_8_32_6), .Cin(s_9_32_6), .S(s_5_32_5), .Cout(s_11_33_5));
    FA FA168 (.A(s_10_32_6), .B(s_11_32_6), .Cin(s_12_32_6), .S(s_4_32_5), .Cout(s_10_33_5));
    FA FA169 (.A(s_13_32_6), .B(s_14_32_6), .Cin(s_15_32_6), .S(s_3_32_5), .Cout(s_9_33_5));
    FA FA170 (.A(s_16_32_6), .B(s_17_32_6), .Cin(s_18_32_6), .S(s_2_32_5), .Cout(s_8_33_5));
    assign s_1_32_5 = s_19_32_6;
    // total 6 half adders and 93 full adders
    // d_6 = 13 done

    assign s_1_1_4 = s_1_1_5;
    assign s_2_2_4 = s_1_2_5;
    assign s_1_2_4 = s_2_2_5;
    assign s_3_3_4 = s_1_3_5;
    assign s_2_3_4 = s_2_3_5;
    assign s_1_3_4 = s_3_3_5;
    assign s_4_4_4 = s_1_4_5;
    assign s_3_4_4 = s_2_4_5;
    assign s_2_4_4 = s_3_4_5;
    assign s_1_4_4 = s_4_4_5;
    assign s_5_5_4 = s_1_5_5;
    assign s_4_5_4 = s_2_5_5;
    assign s_3_5_4 = s_3_5_5;
    assign s_2_5_4 = s_4_5_5;
    assign s_1_5_4 = s_5_5_5;
    assign s_6_6_4 = s_1_6_5;
    assign s_5_6_4 = s_2_6_5;
    assign s_4_6_4 = s_3_6_5;
    assign s_3_6_4 = s_4_6_5;
    assign s_2_6_4 = s_5_6_5;
    assign s_1_6_4 = s_6_6_5;
    assign s_7_7_4 = s_1_7_5;
    assign s_6_7_4 = s_2_7_5;
    assign s_5_7_4 = s_3_7_5;
    assign s_4_7_4 = s_4_7_5;
    assign s_3_7_4 = s_5_7_5;
    assign s_2_7_4 = s_6_7_5;
    assign s_1_7_4 = s_7_7_5;
    assign s_8_8_4 = s_1_8_5;
    assign s_7_8_4 = s_2_8_5;
    assign s_6_8_4 = s_3_8_5;
    assign s_5_8_4 = s_4_8_5;
    assign s_4_8_4 = s_5_8_5;
    assign s_3_8_4 = s_6_8_5;
    assign s_2_8_4 = s_7_8_5;
    assign s_1_8_4 = s_8_8_5;
    assign s_9_9_4 = s_1_9_5;
    assign s_8_9_4 = s_2_9_5;
    assign s_7_9_4 = s_3_9_5;
    assign s_6_9_4 = s_4_9_5;
    assign s_5_9_4 = s_5_9_5;
    assign s_4_9_4 = s_6_9_5;
    assign s_3_9_4 = s_7_9_5;
    assign s_2_9_4 = s_8_9_5;
    assign s_1_9_4 = s_9_9_5;
    HA HA19 (.A(s_1_10_5), .B(s_2_10_5), .S(s_9_10_4), .C(s_9_11_4));
    assign s_8_10_4 = s_3_10_5;
    assign s_7_10_4 = s_4_10_5;
    assign s_6_10_4 = s_5_10_5;
    assign s_5_10_4 = s_6_10_5;
    assign s_4_10_4 = s_7_10_5;
    assign s_3_10_4 = s_8_10_5;
    assign s_2_10_4 = s_9_10_5;
    assign s_1_10_4 = s_10_10_5;
    FA FA171 (.A(s_1_11_5), .B(s_2_11_5), .Cin(s_3_11_5), .S(s_8_11_4), .Cout(s_9_12_4));
    HA HA20 (.A(s_4_11_5), .B(s_5_11_5), .S(s_7_11_4), .C(s_8_12_4));
    assign s_6_11_4 = s_6_11_5;
    assign s_5_11_4 = s_7_11_5;
    assign s_4_11_4 = s_8_11_5;
    assign s_3_11_4 = s_9_11_5;
    assign s_2_11_4 = s_10_11_5;
    assign s_1_11_4 = s_11_11_5;
    FA FA172 (.A(s_1_12_5), .B(s_2_12_5), .Cin(s_3_12_5), .S(s_7_12_4), .Cout(s_9_13_4));
    FA FA173 (.A(s_4_12_5), .B(s_5_12_5), .Cin(s_6_12_5), .S(s_6_12_4), .Cout(s_8_13_4));
    HA HA21 (.A(s_7_12_5), .B(s_8_12_5), .S(s_5_12_4), .C(s_7_13_4));
    assign s_4_12_4 = s_9_12_5;
    assign s_3_12_4 = s_10_12_5;
    assign s_2_12_4 = s_11_12_5;
    assign s_1_12_4 = s_12_12_5;
    FA FA174 (.A(s_1_13_5), .B(s_2_13_5), .Cin(s_3_13_5), .S(s_6_13_4), .Cout(s_9_14_4));
    FA FA175 (.A(s_4_13_5), .B(s_5_13_5), .Cin(s_6_13_5), .S(s_5_13_4), .Cout(s_8_14_4));
    FA FA176 (.A(s_7_13_5), .B(s_8_13_5), .Cin(s_9_13_5), .S(s_4_13_4), .Cout(s_7_14_4));
    HA HA22 (.A(s_10_13_5), .B(s_11_13_5), .S(s_3_13_4), .C(s_6_14_4));
    assign s_2_13_4 = s_12_13_5;
    assign s_1_13_4 = s_13_13_5;
    FA FA177 (.A(s_1_14_5), .B(s_2_14_5), .Cin(s_3_14_5), .S(s_5_14_4), .Cout(s_9_15_4));
    FA FA178 (.A(s_4_14_5), .B(s_5_14_5), .Cin(s_6_14_5), .S(s_4_14_4), .Cout(s_8_15_4));
    FA FA179 (.A(s_7_14_5), .B(s_8_14_5), .Cin(s_9_14_5), .S(s_3_14_4), .Cout(s_7_15_4));
    FA FA180 (.A(s_10_14_5), .B(s_11_14_5), .Cin(s_12_14_5), .S(s_2_14_4), .Cout(s_6_15_4));
    assign s_1_14_4 = s_13_14_5;
    FA FA181 (.A(s_1_15_5), .B(s_2_15_5), .Cin(s_3_15_5), .S(s_5_15_4), .Cout(s_9_16_4));
    FA FA182 (.A(s_4_15_5), .B(s_5_15_5), .Cin(s_6_15_5), .S(s_4_15_4), .Cout(s_8_16_4));
    FA FA183 (.A(s_7_15_5), .B(s_8_15_5), .Cin(s_9_15_5), .S(s_3_15_4), .Cout(s_7_16_4));
    FA FA184 (.A(s_10_15_5), .B(s_11_15_5), .Cin(s_12_15_5), .S(s_2_15_4), .Cout(s_6_16_4));
    assign s_1_15_4 = s_13_15_5;
    FA FA185 (.A(s_1_16_5), .B(s_2_16_5), .Cin(s_3_16_5), .S(s_5_16_4), .Cout(s_9_17_4));
    FA FA186 (.A(s_4_16_5), .B(s_5_16_5), .Cin(s_6_16_5), .S(s_4_16_4), .Cout(s_8_17_4));
    FA FA187 (.A(s_7_16_5), .B(s_8_16_5), .Cin(s_9_16_5), .S(s_3_16_4), .Cout(s_7_17_4));
    FA FA188 (.A(s_10_16_5), .B(s_11_16_5), .Cin(s_12_16_5), .S(s_2_16_4), .Cout(s_6_17_4));
    assign s_1_16_4 = s_13_16_5;
    FA FA189 (.A(s_1_17_5), .B(s_2_17_5), .Cin(s_3_17_5), .S(s_5_17_4), .Cout(s_9_18_4));
    FA FA190 (.A(s_4_17_5), .B(s_5_17_5), .Cin(s_6_17_5), .S(s_4_17_4), .Cout(s_8_18_4));
    FA FA191 (.A(s_7_17_5), .B(s_8_17_5), .Cin(s_9_17_5), .S(s_3_17_4), .Cout(s_7_18_4));
    FA FA192 (.A(s_10_17_5), .B(s_11_17_5), .Cin(s_12_17_5), .S(s_2_17_4), .Cout(s_6_18_4));
    assign s_1_17_4 = s_13_17_5;
    FA FA193 (.A(s_1_18_5), .B(s_2_18_5), .Cin(s_3_18_5), .S(s_5_18_4), .Cout(s_9_19_4));
    FA FA194 (.A(s_4_18_5), .B(s_5_18_5), .Cin(s_6_18_5), .S(s_4_18_4), .Cout(s_8_19_4));
    FA FA195 (.A(s_7_18_5), .B(s_8_18_5), .Cin(s_9_18_5), .S(s_3_18_4), .Cout(s_7_19_4));
    FA FA196 (.A(s_10_18_5), .B(s_11_18_5), .Cin(s_12_18_5), .S(s_2_18_4), .Cout(s_6_19_4));
    assign s_1_18_4 = s_13_18_5;
    FA FA197 (.A(s_1_19_5), .B(s_2_19_5), .Cin(s_3_19_5), .S(s_5_19_4), .Cout(s_9_20_4));
    FA FA198 (.A(s_4_19_5), .B(s_5_19_5), .Cin(s_6_19_5), .S(s_4_19_4), .Cout(s_8_20_4));
    FA FA199 (.A(s_7_19_5), .B(s_8_19_5), .Cin(s_9_19_5), .S(s_3_19_4), .Cout(s_7_20_4));
    FA FA200 (.A(s_10_19_5), .B(s_11_19_5), .Cin(s_12_19_5), .S(s_2_19_4), .Cout(s_6_20_4));
    assign s_1_19_4 = s_13_19_5;
    FA FA201 (.A(s_1_20_5), .B(s_2_20_5), .Cin(s_3_20_5), .S(s_5_20_4), .Cout(s_9_21_4));
    FA FA202 (.A(s_4_20_5), .B(s_5_20_5), .Cin(s_6_20_5), .S(s_4_20_4), .Cout(s_8_21_4));
    FA FA203 (.A(s_7_20_5), .B(s_8_20_5), .Cin(s_9_20_5), .S(s_3_20_4), .Cout(s_7_21_4));
    FA FA204 (.A(s_10_20_5), .B(s_11_20_5), .Cin(s_12_20_5), .S(s_2_20_4), .Cout(s_6_21_4));
    assign s_1_20_4 = s_13_20_5;
    FA FA205 (.A(s_1_21_5), .B(s_2_21_5), .Cin(s_3_21_5), .S(s_5_21_4), .Cout(s_9_22_4));
    FA FA206 (.A(s_4_21_5), .B(s_5_21_5), .Cin(s_6_21_5), .S(s_4_21_4), .Cout(s_8_22_4));
    FA FA207 (.A(s_7_21_5), .B(s_8_21_5), .Cin(s_9_21_5), .S(s_3_21_4), .Cout(s_7_22_4));
    FA FA208 (.A(s_10_21_5), .B(s_11_21_5), .Cin(s_12_21_5), .S(s_2_21_4), .Cout(s_6_22_4));
    assign s_1_21_4 = s_13_21_5;
    FA FA209 (.A(s_1_22_5), .B(s_2_22_5), .Cin(s_3_22_5), .S(s_5_22_4), .Cout(s_9_23_4));
    FA FA210 (.A(s_4_22_5), .B(s_5_22_5), .Cin(s_6_22_5), .S(s_4_22_4), .Cout(s_8_23_4));
    FA FA211 (.A(s_7_22_5), .B(s_8_22_5), .Cin(s_9_22_5), .S(s_3_22_4), .Cout(s_7_23_4));
    FA FA212 (.A(s_10_22_5), .B(s_11_22_5), .Cin(s_12_22_5), .S(s_2_22_4), .Cout(s_6_23_4));
    assign s_1_22_4 = s_13_22_5;
    FA FA213 (.A(s_1_23_5), .B(s_2_23_5), .Cin(s_3_23_5), .S(s_5_23_4), .Cout(s_9_24_4));
    FA FA214 (.A(s_4_23_5), .B(s_5_23_5), .Cin(s_6_23_5), .S(s_4_23_4), .Cout(s_8_24_4));
    FA FA215 (.A(s_7_23_5), .B(s_8_23_5), .Cin(s_9_23_5), .S(s_3_23_4), .Cout(s_7_24_4));
    FA FA216 (.A(s_10_23_5), .B(s_11_23_5), .Cin(s_12_23_5), .S(s_2_23_4), .Cout(s_6_24_4));
    assign s_1_23_4 = s_13_23_5;
    FA FA217 (.A(s_1_24_5), .B(s_2_24_5), .Cin(s_3_24_5), .S(s_5_24_4), .Cout(s_9_25_4));
    FA FA218 (.A(s_4_24_5), .B(s_5_24_5), .Cin(s_6_24_5), .S(s_4_24_4), .Cout(s_8_25_4));
    FA FA219 (.A(s_7_24_5), .B(s_8_24_5), .Cin(s_9_24_5), .S(s_3_24_4), .Cout(s_7_25_4));
    FA FA220 (.A(s_10_24_5), .B(s_11_24_5), .Cin(s_12_24_5), .S(s_2_24_4), .Cout(s_6_25_4));
    assign s_1_24_4 = s_13_24_5;
    FA FA221 (.A(s_1_25_5), .B(s_2_25_5), .Cin(s_3_25_5), .S(s_5_25_4), .Cout(s_9_26_4));
    FA FA222 (.A(s_4_25_5), .B(s_5_25_5), .Cin(s_6_25_5), .S(s_4_25_4), .Cout(s_8_26_4));
    FA FA223 (.A(s_7_25_5), .B(s_8_25_5), .Cin(s_9_25_5), .S(s_3_25_4), .Cout(s_7_26_4));
    FA FA224 (.A(s_10_25_5), .B(s_11_25_5), .Cin(s_12_25_5), .S(s_2_25_4), .Cout(s_6_26_4));
    assign s_1_25_4 = s_13_25_5;
    FA FA225 (.A(s_1_26_5), .B(s_2_26_5), .Cin(s_3_26_5), .S(s_5_26_4), .Cout(s_9_27_4));
    FA FA226 (.A(s_4_26_5), .B(s_5_26_5), .Cin(s_6_26_5), .S(s_4_26_4), .Cout(s_8_27_4));
    FA FA227 (.A(s_7_26_5), .B(s_8_26_5), .Cin(s_9_26_5), .S(s_3_26_4), .Cout(s_7_27_4));
    FA FA228 (.A(s_10_26_5), .B(s_11_26_5), .Cin(s_12_26_5), .S(s_2_26_4), .Cout(s_6_27_4));
    assign s_1_26_4 = s_13_26_5;
    FA FA229 (.A(s_1_27_5), .B(s_2_27_5), .Cin(s_3_27_5), .S(s_5_27_4), .Cout(s_9_28_4));
    FA FA230 (.A(s_4_27_5), .B(s_5_27_5), .Cin(s_6_27_5), .S(s_4_27_4), .Cout(s_8_28_4));
    FA FA231 (.A(s_7_27_5), .B(s_8_27_5), .Cin(s_9_27_5), .S(s_3_27_4), .Cout(s_7_28_4));
    FA FA232 (.A(s_10_27_5), .B(s_11_27_5), .Cin(s_12_27_5), .S(s_2_27_4), .Cout(s_6_28_4));
    assign s_1_27_4 = s_13_27_5;
    FA FA233 (.A(s_1_28_5), .B(s_2_28_5), .Cin(s_3_28_5), .S(s_5_28_4), .Cout(s_9_29_4));
    FA FA234 (.A(s_4_28_5), .B(s_5_28_5), .Cin(s_6_28_5), .S(s_4_28_4), .Cout(s_8_29_4));
    FA FA235 (.A(s_7_28_5), .B(s_8_28_5), .Cin(s_9_28_5), .S(s_3_28_4), .Cout(s_7_29_4));
    FA FA236 (.A(s_10_28_5), .B(s_11_28_5), .Cin(s_12_28_5), .S(s_2_28_4), .Cout(s_6_29_4));
    assign s_1_28_4 = s_13_28_5;
    FA FA237 (.A(s_1_29_5), .B(s_2_29_5), .Cin(s_3_29_5), .S(s_5_29_4), .Cout(s_9_30_4));
    FA FA238 (.A(s_4_29_5), .B(s_5_29_5), .Cin(s_6_29_5), .S(s_4_29_4), .Cout(s_8_30_4));
    FA FA239 (.A(s_7_29_5), .B(s_8_29_5), .Cin(s_9_29_5), .S(s_3_29_4), .Cout(s_7_30_4));
    FA FA240 (.A(s_10_29_5), .B(s_11_29_5), .Cin(s_12_29_5), .S(s_2_29_4), .Cout(s_6_30_4));
    assign s_1_29_4 = s_13_29_5;
    FA FA241 (.A(s_1_30_5), .B(s_2_30_5), .Cin(s_3_30_5), .S(s_5_30_4), .Cout(s_9_31_4));
    FA FA242 (.A(s_4_30_5), .B(s_5_30_5), .Cin(s_6_30_5), .S(s_4_30_4), .Cout(s_8_31_4));
    FA FA243 (.A(s_7_30_5), .B(s_8_30_5), .Cin(s_9_30_5), .S(s_3_30_4), .Cout(s_7_31_4));
    FA FA244 (.A(s_10_30_5), .B(s_11_30_5), .Cin(s_12_30_5), .S(s_2_30_4), .Cout(s_6_31_4));
    assign s_1_30_4 = s_13_30_5;
    FA FA245 (.A(s_1_31_5), .B(s_2_31_5), .Cin(s_3_31_5), .S(s_5_31_4), .Cout(s_9_32_4));
    FA FA246 (.A(s_4_31_5), .B(s_5_31_5), .Cin(s_6_31_5), .S(s_4_31_4), .Cout(s_8_32_4));
    FA FA247 (.A(s_7_31_5), .B(s_8_31_5), .Cin(s_9_31_5), .S(s_3_31_4), .Cout(s_7_32_4));
    FA FA248 (.A(s_10_31_5), .B(s_11_31_5), .Cin(s_12_31_5), .S(s_2_31_4), .Cout(s_6_32_4));
    assign s_1_31_4 = s_13_31_5;
    FA FA249 (.A(s_1_32_5), .B(s_2_32_5), .Cin(s_3_32_5), .S(s_5_32_4), .Cout(s_9_33_4));
    FA FA250 (.A(s_4_32_5), .B(s_5_32_5), .Cin(s_6_32_5), .S(s_4_32_4), .Cout(s_8_33_4));
    FA FA251 (.A(s_7_32_5), .B(s_8_32_5), .Cin(s_9_32_5), .S(s_3_32_4), .Cout(s_7_33_4));
    FA FA252 (.A(s_10_32_5), .B(s_11_32_5), .Cin(s_12_32_5), .S(s_2_32_4), .Cout(s_6_33_4));
    assign s_1_32_4 = s_13_32_5;
    // total 4 half adders and 82 full adders
    // d_5 = 9 done

    assign s_1_1_3 = s_1_1_4;
    assign s_2_2_3 = s_1_2_4;
    assign s_1_2_3 = s_2_2_4;
    assign s_3_3_3 = s_1_3_4;
    assign s_2_3_3 = s_2_3_4;
    assign s_1_3_3 = s_3_3_4;
    assign s_4_4_3 = s_1_4_4;
    assign s_3_4_3 = s_2_4_4;
    assign s_2_4_3 = s_3_4_4;
    assign s_1_4_3 = s_4_4_4;
    assign s_5_5_3 = s_1_5_4;
    assign s_4_5_3 = s_2_5_4;
    assign s_3_5_3 = s_3_5_4;
    assign s_2_5_3 = s_4_5_4;
    assign s_1_5_3 = s_5_5_4;
    assign s_6_6_3 = s_1_6_4;
    assign s_5_6_3 = s_2_6_4;
    assign s_4_6_3 = s_3_6_4;
    assign s_3_6_3 = s_4_6_4;
    assign s_2_6_3 = s_5_6_4;
    assign s_1_6_3 = s_6_6_4;
    HA HA23 (.A(s_1_7_4), .B(s_2_7_4), .S(s_6_7_3), .C(s_6_8_3));
    assign s_5_7_3 = s_3_7_4;
    assign s_4_7_3 = s_4_7_4;
    assign s_3_7_3 = s_5_7_4;
    assign s_2_7_3 = s_6_7_4;
    assign s_1_7_3 = s_7_7_4;
    FA FA253 (.A(s_1_8_4), .B(s_2_8_4), .Cin(s_3_8_4), .S(s_5_8_3), .Cout(s_6_9_3));
    HA HA24 (.A(s_4_8_4), .B(s_5_8_4), .S(s_4_8_3), .C(s_5_9_3));
    assign s_3_8_3 = s_6_8_4;
    assign s_2_8_3 = s_7_8_4;
    assign s_1_8_3 = s_8_8_4;
    FA FA254 (.A(s_1_9_4), .B(s_2_9_4), .Cin(s_3_9_4), .S(s_4_9_3), .Cout(s_6_10_3));
    FA FA255 (.A(s_4_9_4), .B(s_5_9_4), .Cin(s_6_9_4), .S(s_3_9_3), .Cout(s_5_10_3));
    HA HA25 (.A(s_7_9_4), .B(s_8_9_4), .S(s_2_9_3), .C(s_4_10_3));
    assign s_1_9_3 = s_9_9_4;
    FA FA256 (.A(s_1_10_4), .B(s_2_10_4), .Cin(s_3_10_4), .S(s_3_10_3), .Cout(s_6_11_3));
    FA FA257 (.A(s_4_10_4), .B(s_5_10_4), .Cin(s_6_10_4), .S(s_2_10_3), .Cout(s_5_11_3));
    FA FA258 (.A(s_7_10_4), .B(s_8_10_4), .Cin(s_9_10_4), .S(s_1_10_3), .Cout(s_4_11_3));
    FA FA259 (.A(s_1_11_4), .B(s_2_11_4), .Cin(s_3_11_4), .S(s_3_11_3), .Cout(s_6_12_3));
    FA FA260 (.A(s_4_11_4), .B(s_5_11_4), .Cin(s_6_11_4), .S(s_2_11_3), .Cout(s_5_12_3));
    FA FA261 (.A(s_7_11_4), .B(s_8_11_4), .Cin(s_9_11_4), .S(s_1_11_3), .Cout(s_4_12_3));
    FA FA262 (.A(s_1_12_4), .B(s_2_12_4), .Cin(s_3_12_4), .S(s_3_12_3), .Cout(s_6_13_3));
    FA FA263 (.A(s_4_12_4), .B(s_5_12_4), .Cin(s_6_12_4), .S(s_2_12_3), .Cout(s_5_13_3));
    FA FA264 (.A(s_7_12_4), .B(s_8_12_4), .Cin(s_9_12_4), .S(s_1_12_3), .Cout(s_4_13_3));
    FA FA265 (.A(s_1_13_4), .B(s_2_13_4), .Cin(s_3_13_4), .S(s_3_13_3), .Cout(s_6_14_3));
    FA FA266 (.A(s_4_13_4), .B(s_5_13_4), .Cin(s_6_13_4), .S(s_2_13_3), .Cout(s_5_14_3));
    FA FA267 (.A(s_7_13_4), .B(s_8_13_4), .Cin(s_9_13_4), .S(s_1_13_3), .Cout(s_4_14_3));
    FA FA268 (.A(s_1_14_4), .B(s_2_14_4), .Cin(s_3_14_4), .S(s_3_14_3), .Cout(s_6_15_3));
    FA FA269 (.A(s_4_14_4), .B(s_5_14_4), .Cin(s_6_14_4), .S(s_2_14_3), .Cout(s_5_15_3));
    FA FA270 (.A(s_7_14_4), .B(s_8_14_4), .Cin(s_9_14_4), .S(s_1_14_3), .Cout(s_4_15_3));
    FA FA271 (.A(s_1_15_4), .B(s_2_15_4), .Cin(s_3_15_4), .S(s_3_15_3), .Cout(s_6_16_3));
    FA FA272 (.A(s_4_15_4), .B(s_5_15_4), .Cin(s_6_15_4), .S(s_2_15_3), .Cout(s_5_16_3));
    FA FA273 (.A(s_7_15_4), .B(s_8_15_4), .Cin(s_9_15_4), .S(s_1_15_3), .Cout(s_4_16_3));
    FA FA274 (.A(s_1_16_4), .B(s_2_16_4), .Cin(s_3_16_4), .S(s_3_16_3), .Cout(s_6_17_3));
    FA FA275 (.A(s_4_16_4), .B(s_5_16_4), .Cin(s_6_16_4), .S(s_2_16_3), .Cout(s_5_17_3));
    FA FA276 (.A(s_7_16_4), .B(s_8_16_4), .Cin(s_9_16_4), .S(s_1_16_3), .Cout(s_4_17_3));
    FA FA277 (.A(s_1_17_4), .B(s_2_17_4), .Cin(s_3_17_4), .S(s_3_17_3), .Cout(s_6_18_3));
    FA FA278 (.A(s_4_17_4), .B(s_5_17_4), .Cin(s_6_17_4), .S(s_2_17_3), .Cout(s_5_18_3));
    FA FA279 (.A(s_7_17_4), .B(s_8_17_4), .Cin(s_9_17_4), .S(s_1_17_3), .Cout(s_4_18_3));
    FA FA280 (.A(s_1_18_4), .B(s_2_18_4), .Cin(s_3_18_4), .S(s_3_18_3), .Cout(s_6_19_3));
    FA FA281 (.A(s_4_18_4), .B(s_5_18_4), .Cin(s_6_18_4), .S(s_2_18_3), .Cout(s_5_19_3));
    FA FA282 (.A(s_7_18_4), .B(s_8_18_4), .Cin(s_9_18_4), .S(s_1_18_3), .Cout(s_4_19_3));
    FA FA283 (.A(s_1_19_4), .B(s_2_19_4), .Cin(s_3_19_4), .S(s_3_19_3), .Cout(s_6_20_3));
    FA FA284 (.A(s_4_19_4), .B(s_5_19_4), .Cin(s_6_19_4), .S(s_2_19_3), .Cout(s_5_20_3));
    FA FA285 (.A(s_7_19_4), .B(s_8_19_4), .Cin(s_9_19_4), .S(s_1_19_3), .Cout(s_4_20_3));
    FA FA286 (.A(s_1_20_4), .B(s_2_20_4), .Cin(s_3_20_4), .S(s_3_20_3), .Cout(s_6_21_3));
    FA FA287 (.A(s_4_20_4), .B(s_5_20_4), .Cin(s_6_20_4), .S(s_2_20_3), .Cout(s_5_21_3));
    FA FA288 (.A(s_7_20_4), .B(s_8_20_4), .Cin(s_9_20_4), .S(s_1_20_3), .Cout(s_4_21_3));
    FA FA289 (.A(s_1_21_4), .B(s_2_21_4), .Cin(s_3_21_4), .S(s_3_21_3), .Cout(s_6_22_3));
    FA FA290 (.A(s_4_21_4), .B(s_5_21_4), .Cin(s_6_21_4), .S(s_2_21_3), .Cout(s_5_22_3));
    FA FA291 (.A(s_7_21_4), .B(s_8_21_4), .Cin(s_9_21_4), .S(s_1_21_3), .Cout(s_4_22_3));
    FA FA292 (.A(s_1_22_4), .B(s_2_22_4), .Cin(s_3_22_4), .S(s_3_22_3), .Cout(s_6_23_3));
    FA FA293 (.A(s_4_22_4), .B(s_5_22_4), .Cin(s_6_22_4), .S(s_2_22_3), .Cout(s_5_23_3));
    FA FA294 (.A(s_7_22_4), .B(s_8_22_4), .Cin(s_9_22_4), .S(s_1_22_3), .Cout(s_4_23_3));
    FA FA295 (.A(s_1_23_4), .B(s_2_23_4), .Cin(s_3_23_4), .S(s_3_23_3), .Cout(s_6_24_3));
    FA FA296 (.A(s_4_23_4), .B(s_5_23_4), .Cin(s_6_23_4), .S(s_2_23_3), .Cout(s_5_24_3));
    FA FA297 (.A(s_7_23_4), .B(s_8_23_4), .Cin(s_9_23_4), .S(s_1_23_3), .Cout(s_4_24_3));
    FA FA298 (.A(s_1_24_4), .B(s_2_24_4), .Cin(s_3_24_4), .S(s_3_24_3), .Cout(s_6_25_3));
    FA FA299 (.A(s_4_24_4), .B(s_5_24_4), .Cin(s_6_24_4), .S(s_2_24_3), .Cout(s_5_25_3));
    FA FA300 (.A(s_7_24_4), .B(s_8_24_4), .Cin(s_9_24_4), .S(s_1_24_3), .Cout(s_4_25_3));
    FA FA301 (.A(s_1_25_4), .B(s_2_25_4), .Cin(s_3_25_4), .S(s_3_25_3), .Cout(s_6_26_3));
    FA FA302 (.A(s_4_25_4), .B(s_5_25_4), .Cin(s_6_25_4), .S(s_2_25_3), .Cout(s_5_26_3));
    FA FA303 (.A(s_7_25_4), .B(s_8_25_4), .Cin(s_9_25_4), .S(s_1_25_3), .Cout(s_4_26_3));
    FA FA304 (.A(s_1_26_4), .B(s_2_26_4), .Cin(s_3_26_4), .S(s_3_26_3), .Cout(s_6_27_3));
    FA FA305 (.A(s_4_26_4), .B(s_5_26_4), .Cin(s_6_26_4), .S(s_2_26_3), .Cout(s_5_27_3));
    FA FA306 (.A(s_7_26_4), .B(s_8_26_4), .Cin(s_9_26_4), .S(s_1_26_3), .Cout(s_4_27_3));
    FA FA307 (.A(s_1_27_4), .B(s_2_27_4), .Cin(s_3_27_4), .S(s_3_27_3), .Cout(s_6_28_3));
    FA FA308 (.A(s_4_27_4), .B(s_5_27_4), .Cin(s_6_27_4), .S(s_2_27_3), .Cout(s_5_28_3));
    FA FA309 (.A(s_7_27_4), .B(s_8_27_4), .Cin(s_9_27_4), .S(s_1_27_3), .Cout(s_4_28_3));
    FA FA310 (.A(s_1_28_4), .B(s_2_28_4), .Cin(s_3_28_4), .S(s_3_28_3), .Cout(s_6_29_3));
    FA FA311 (.A(s_4_28_4), .B(s_5_28_4), .Cin(s_6_28_4), .S(s_2_28_3), .Cout(s_5_29_3));
    FA FA312 (.A(s_7_28_4), .B(s_8_28_4), .Cin(s_9_28_4), .S(s_1_28_3), .Cout(s_4_29_3));
    FA FA313 (.A(s_1_29_4), .B(s_2_29_4), .Cin(s_3_29_4), .S(s_3_29_3), .Cout(s_6_30_3));
    FA FA314 (.A(s_4_29_4), .B(s_5_29_4), .Cin(s_6_29_4), .S(s_2_29_3), .Cout(s_5_30_3));
    FA FA315 (.A(s_7_29_4), .B(s_8_29_4), .Cin(s_9_29_4), .S(s_1_29_3), .Cout(s_4_30_3));
    FA FA316 (.A(s_1_30_4), .B(s_2_30_4), .Cin(s_3_30_4), .S(s_3_30_3), .Cout(s_6_31_3));
    FA FA317 (.A(s_4_30_4), .B(s_5_30_4), .Cin(s_6_30_4), .S(s_2_30_3), .Cout(s_5_31_3));
    FA FA318 (.A(s_7_30_4), .B(s_8_30_4), .Cin(s_9_30_4), .S(s_1_30_3), .Cout(s_4_31_3));
    FA FA319 (.A(s_1_31_4), .B(s_2_31_4), .Cin(s_3_31_4), .S(s_3_31_3), .Cout(s_6_32_3));
    FA FA320 (.A(s_4_31_4), .B(s_5_31_4), .Cin(s_6_31_4), .S(s_2_31_3), .Cout(s_5_32_3));
    FA FA321 (.A(s_7_31_4), .B(s_8_31_4), .Cin(s_9_31_4), .S(s_1_31_3), .Cout(s_4_32_3));
    FA FA322 (.A(s_1_32_4), .B(s_2_32_4), .Cin(s_3_32_4), .S(s_3_32_3), .Cout(s_6_33_3));
    FA FA323 (.A(s_4_32_4), .B(s_5_32_4), .Cin(s_6_32_4), .S(s_2_32_3), .Cout(s_5_33_3));
    FA FA324 (.A(s_7_32_4), .B(s_8_32_4), .Cin(s_9_32_4), .S(s_1_32_3), .Cout(s_4_33_3));
    // total 3 half adders and 72 full adders
    // d_4 = 6 done

    assign s_1_1_2 = s_1_1_3;
    assign s_2_2_2 = s_1_2_3;
    assign s_1_2_2 = s_2_2_3;
    assign s_3_3_2 = s_1_3_3;
    assign s_2_3_2 = s_2_3_3;
    assign s_1_3_2 = s_3_3_3;
    assign s_4_4_2 = s_1_4_3;
    assign s_3_4_2 = s_2_4_3;
    assign s_2_4_2 = s_3_4_3;
    assign s_1_4_2 = s_4_4_3;
    HA HA26 (.A(s_1_5_3), .B(s_2_5_3), .S(s_4_5_2), .C(s_4_6_2));
    assign s_3_5_2 = s_3_5_3;
    assign s_2_5_2 = s_4_5_3;
    assign s_1_5_2 = s_5_5_3;
    FA FA325 (.A(s_1_6_3), .B(s_2_6_3), .Cin(s_3_6_3), .S(s_3_6_2), .Cout(s_4_7_2));
    HA HA27 (.A(s_4_6_3), .B(s_5_6_3), .S(s_2_6_2), .C(s_3_7_2));
    assign s_1_6_2 = s_6_6_3;
    FA FA326 (.A(s_1_7_3), .B(s_2_7_3), .Cin(s_3_7_3), .S(s_2_7_2), .Cout(s_4_8_2));
    FA FA327 (.A(s_4_7_3), .B(s_5_7_3), .Cin(s_6_7_3), .S(s_1_7_2), .Cout(s_3_8_2));
    FA FA328 (.A(s_1_8_3), .B(s_2_8_3), .Cin(s_3_8_3), .S(s_2_8_2), .Cout(s_4_9_2));
    FA FA329 (.A(s_4_8_3), .B(s_5_8_3), .Cin(s_6_8_3), .S(s_1_8_2), .Cout(s_3_9_2));
    FA FA330 (.A(s_1_9_3), .B(s_2_9_3), .Cin(s_3_9_3), .S(s_2_9_2), .Cout(s_4_10_2));
    FA FA331 (.A(s_4_9_3), .B(s_5_9_3), .Cin(s_6_9_3), .S(s_1_9_2), .Cout(s_3_10_2));
    FA FA332 (.A(s_1_10_3), .B(s_2_10_3), .Cin(s_3_10_3), .S(s_2_10_2), .Cout(s_4_11_2));
    FA FA333 (.A(s_4_10_3), .B(s_5_10_3), .Cin(s_6_10_3), .S(s_1_10_2), .Cout(s_3_11_2));
    FA FA334 (.A(s_1_11_3), .B(s_2_11_3), .Cin(s_3_11_3), .S(s_2_11_2), .Cout(s_4_12_2));
    FA FA335 (.A(s_4_11_3), .B(s_5_11_3), .Cin(s_6_11_3), .S(s_1_11_2), .Cout(s_3_12_2));
    FA FA336 (.A(s_1_12_3), .B(s_2_12_3), .Cin(s_3_12_3), .S(s_2_12_2), .Cout(s_4_13_2));
    FA FA337 (.A(s_4_12_3), .B(s_5_12_3), .Cin(s_6_12_3), .S(s_1_12_2), .Cout(s_3_13_2));
    FA FA338 (.A(s_1_13_3), .B(s_2_13_3), .Cin(s_3_13_3), .S(s_2_13_2), .Cout(s_4_14_2));
    FA FA339 (.A(s_4_13_3), .B(s_5_13_3), .Cin(s_6_13_3), .S(s_1_13_2), .Cout(s_3_14_2));
    FA FA340 (.A(s_1_14_3), .B(s_2_14_3), .Cin(s_3_14_3), .S(s_2_14_2), .Cout(s_4_15_2));
    FA FA341 (.A(s_4_14_3), .B(s_5_14_3), .Cin(s_6_14_3), .S(s_1_14_2), .Cout(s_3_15_2));
    FA FA342 (.A(s_1_15_3), .B(s_2_15_3), .Cin(s_3_15_3), .S(s_2_15_2), .Cout(s_4_16_2));
    FA FA343 (.A(s_4_15_3), .B(s_5_15_3), .Cin(s_6_15_3), .S(s_1_15_2), .Cout(s_3_16_2));
    FA FA344 (.A(s_1_16_3), .B(s_2_16_3), .Cin(s_3_16_3), .S(s_2_16_2), .Cout(s_4_17_2));
    FA FA345 (.A(s_4_16_3), .B(s_5_16_3), .Cin(s_6_16_3), .S(s_1_16_2), .Cout(s_3_17_2));
    FA FA346 (.A(s_1_17_3), .B(s_2_17_3), .Cin(s_3_17_3), .S(s_2_17_2), .Cout(s_4_18_2));
    FA FA347 (.A(s_4_17_3), .B(s_5_17_3), .Cin(s_6_17_3), .S(s_1_17_2), .Cout(s_3_18_2));
    FA FA348 (.A(s_1_18_3), .B(s_2_18_3), .Cin(s_3_18_3), .S(s_2_18_2), .Cout(s_4_19_2));
    FA FA349 (.A(s_4_18_3), .B(s_5_18_3), .Cin(s_6_18_3), .S(s_1_18_2), .Cout(s_3_19_2));
    FA FA350 (.A(s_1_19_3), .B(s_2_19_3), .Cin(s_3_19_3), .S(s_2_19_2), .Cout(s_4_20_2));
    FA FA351 (.A(s_4_19_3), .B(s_5_19_3), .Cin(s_6_19_3), .S(s_1_19_2), .Cout(s_3_20_2));
    FA FA352 (.A(s_1_20_3), .B(s_2_20_3), .Cin(s_3_20_3), .S(s_2_20_2), .Cout(s_4_21_2));
    FA FA353 (.A(s_4_20_3), .B(s_5_20_3), .Cin(s_6_20_3), .S(s_1_20_2), .Cout(s_3_21_2));
    FA FA354 (.A(s_1_21_3), .B(s_2_21_3), .Cin(s_3_21_3), .S(s_2_21_2), .Cout(s_4_22_2));
    FA FA355 (.A(s_4_21_3), .B(s_5_21_3), .Cin(s_6_21_3), .S(s_1_21_2), .Cout(s_3_22_2));
    FA FA356 (.A(s_1_22_3), .B(s_2_22_3), .Cin(s_3_22_3), .S(s_2_22_2), .Cout(s_4_23_2));
    FA FA357 (.A(s_4_22_3), .B(s_5_22_3), .Cin(s_6_22_3), .S(s_1_22_2), .Cout(s_3_23_2));
    FA FA358 (.A(s_1_23_3), .B(s_2_23_3), .Cin(s_3_23_3), .S(s_2_23_2), .Cout(s_4_24_2));
    FA FA359 (.A(s_4_23_3), .B(s_5_23_3), .Cin(s_6_23_3), .S(s_1_23_2), .Cout(s_3_24_2));
    FA FA360 (.A(s_1_24_3), .B(s_2_24_3), .Cin(s_3_24_3), .S(s_2_24_2), .Cout(s_4_25_2));
    FA FA361 (.A(s_4_24_3), .B(s_5_24_3), .Cin(s_6_24_3), .S(s_1_24_2), .Cout(s_3_25_2));
    FA FA362 (.A(s_1_25_3), .B(s_2_25_3), .Cin(s_3_25_3), .S(s_2_25_2), .Cout(s_4_26_2));
    FA FA363 (.A(s_4_25_3), .B(s_5_25_3), .Cin(s_6_25_3), .S(s_1_25_2), .Cout(s_3_26_2));
    FA FA364 (.A(s_1_26_3), .B(s_2_26_3), .Cin(s_3_26_3), .S(s_2_26_2), .Cout(s_4_27_2));
    FA FA365 (.A(s_4_26_3), .B(s_5_26_3), .Cin(s_6_26_3), .S(s_1_26_2), .Cout(s_3_27_2));
    FA FA366 (.A(s_1_27_3), .B(s_2_27_3), .Cin(s_3_27_3), .S(s_2_27_2), .Cout(s_4_28_2));
    FA FA367 (.A(s_4_27_3), .B(s_5_27_3), .Cin(s_6_27_3), .S(s_1_27_2), .Cout(s_3_28_2));
    FA FA368 (.A(s_1_28_3), .B(s_2_28_3), .Cin(s_3_28_3), .S(s_2_28_2), .Cout(s_4_29_2));
    FA FA369 (.A(s_4_28_3), .B(s_5_28_3), .Cin(s_6_28_3), .S(s_1_28_2), .Cout(s_3_29_2));
    FA FA370 (.A(s_1_29_3), .B(s_2_29_3), .Cin(s_3_29_3), .S(s_2_29_2), .Cout(s_4_30_2));
    FA FA371 (.A(s_4_29_3), .B(s_5_29_3), .Cin(s_6_29_3), .S(s_1_29_2), .Cout(s_3_30_2));
    FA FA372 (.A(s_1_30_3), .B(s_2_30_3), .Cin(s_3_30_3), .S(s_2_30_2), .Cout(s_4_31_2));
    FA FA373 (.A(s_4_30_3), .B(s_5_30_3), .Cin(s_6_30_3), .S(s_1_30_2), .Cout(s_3_31_2));
    FA FA374 (.A(s_1_31_3), .B(s_2_31_3), .Cin(s_3_31_3), .S(s_2_31_2), .Cout(s_4_32_2));
    FA FA375 (.A(s_4_31_3), .B(s_5_31_3), .Cin(s_6_31_3), .S(s_1_31_2), .Cout(s_3_32_2));
    FA FA376 (.A(s_1_32_3), .B(s_2_32_3), .Cin(s_3_32_3), .S(s_2_32_2), .Cout(s_4_33_2));
    FA FA377 (.A(s_4_32_3), .B(s_5_32_3), .Cin(s_6_32_3), .S(s_1_32_2), .Cout(s_3_33_2));
    // total 2 half adders and 53 full adders
    // d_3 = 4 done

    assign s_1_1_1 = s_1_1_2;
    assign s_2_2_1 = s_1_2_2;
    assign s_1_2_1 = s_2_2_2;
    assign s_3_3_1 = s_1_3_2;
    assign s_2_3_1 = s_2_3_2;
    assign s_1_3_1 = s_3_3_2;
    HA HA28 (.A(s_1_4_2), .B(s_2_4_2), .S(s_3_4_1), .C(s_3_5_1));
    assign s_2_4_1 = s_3_4_2;
    assign s_1_4_1 = s_4_4_2;
    FA FA378 (.A(s_1_5_2), .B(s_2_5_2), .Cin(s_3_5_2), .S(s_2_5_1), .Cout(s_3_6_1));
    assign s_1_5_1 = s_4_5_2;
    FA FA379 (.A(s_1_6_2), .B(s_2_6_2), .Cin(s_3_6_2), .S(s_2_6_1), .Cout(s_3_7_1));
    assign s_1_6_1 = s_4_6_2;
    FA FA380 (.A(s_1_7_2), .B(s_2_7_2), .Cin(s_3_7_2), .S(s_2_7_1), .Cout(s_3_8_1));
    assign s_1_7_1 = s_4_7_2;
    FA FA381 (.A(s_1_8_2), .B(s_2_8_2), .Cin(s_3_8_2), .S(s_2_8_1), .Cout(s_3_9_1));
    assign s_1_8_1 = s_4_8_2;
    FA FA382 (.A(s_1_9_2), .B(s_2_9_2), .Cin(s_3_9_2), .S(s_2_9_1), .Cout(s_3_10_1));
    assign s_1_9_1 = s_4_9_2;
    FA FA383 (.A(s_1_10_2), .B(s_2_10_2), .Cin(s_3_10_2), .S(s_2_10_1), .Cout(s_3_11_1));
    assign s_1_10_1 = s_4_10_2;
    FA FA384 (.A(s_1_11_2), .B(s_2_11_2), .Cin(s_3_11_2), .S(s_2_11_1), .Cout(s_3_12_1));
    assign s_1_11_1 = s_4_11_2;
    FA FA385 (.A(s_1_12_2), .B(s_2_12_2), .Cin(s_3_12_2), .S(s_2_12_1), .Cout(s_3_13_1));
    assign s_1_12_1 = s_4_12_2;
    FA FA386 (.A(s_1_13_2), .B(s_2_13_2), .Cin(s_3_13_2), .S(s_2_13_1), .Cout(s_3_14_1));
    assign s_1_13_1 = s_4_13_2;
    FA FA387 (.A(s_1_14_2), .B(s_2_14_2), .Cin(s_3_14_2), .S(s_2_14_1), .Cout(s_3_15_1));
    assign s_1_14_1 = s_4_14_2;
    FA FA388 (.A(s_1_15_2), .B(s_2_15_2), .Cin(s_3_15_2), .S(s_2_15_1), .Cout(s_3_16_1));
    assign s_1_15_1 = s_4_15_2;
    FA FA389 (.A(s_1_16_2), .B(s_2_16_2), .Cin(s_3_16_2), .S(s_2_16_1), .Cout(s_3_17_1));
    assign s_1_16_1 = s_4_16_2;
    FA FA390 (.A(s_1_17_2), .B(s_2_17_2), .Cin(s_3_17_2), .S(s_2_17_1), .Cout(s_3_18_1));
    assign s_1_17_1 = s_4_17_2;
    FA FA391 (.A(s_1_18_2), .B(s_2_18_2), .Cin(s_3_18_2), .S(s_2_18_1), .Cout(s_3_19_1));
    assign s_1_18_1 = s_4_18_2;
    FA FA392 (.A(s_1_19_2), .B(s_2_19_2), .Cin(s_3_19_2), .S(s_2_19_1), .Cout(s_3_20_1));
    assign s_1_19_1 = s_4_19_2;
    FA FA393 (.A(s_1_20_2), .B(s_2_20_2), .Cin(s_3_20_2), .S(s_2_20_1), .Cout(s_3_21_1));
    assign s_1_20_1 = s_4_20_2;
    FA FA394 (.A(s_1_21_2), .B(s_2_21_2), .Cin(s_3_21_2), .S(s_2_21_1), .Cout(s_3_22_1));
    assign s_1_21_1 = s_4_21_2;
    FA FA395 (.A(s_1_22_2), .B(s_2_22_2), .Cin(s_3_22_2), .S(s_2_22_1), .Cout(s_3_23_1));
    assign s_1_22_1 = s_4_22_2;
    FA FA396 (.A(s_1_23_2), .B(s_2_23_2), .Cin(s_3_23_2), .S(s_2_23_1), .Cout(s_3_24_1));
    assign s_1_23_1 = s_4_23_2;
    FA FA397 (.A(s_1_24_2), .B(s_2_24_2), .Cin(s_3_24_2), .S(s_2_24_1), .Cout(s_3_25_1));
    assign s_1_24_1 = s_4_24_2;
    FA FA398 (.A(s_1_25_2), .B(s_2_25_2), .Cin(s_3_25_2), .S(s_2_25_1), .Cout(s_3_26_1));
    assign s_1_25_1 = s_4_25_2;
    FA FA399 (.A(s_1_26_2), .B(s_2_26_2), .Cin(s_3_26_2), .S(s_2_26_1), .Cout(s_3_27_1));
    assign s_1_26_1 = s_4_26_2;
    FA FA400 (.A(s_1_27_2), .B(s_2_27_2), .Cin(s_3_27_2), .S(s_2_27_1), .Cout(s_3_28_1));
    assign s_1_27_1 = s_4_27_2;
    FA FA401 (.A(s_1_28_2), .B(s_2_28_2), .Cin(s_3_28_2), .S(s_2_28_1), .Cout(s_3_29_1));
    assign s_1_28_1 = s_4_28_2;
    FA FA402 (.A(s_1_29_2), .B(s_2_29_2), .Cin(s_3_29_2), .S(s_2_29_1), .Cout(s_3_30_1));
    assign s_1_29_1 = s_4_29_2;
    FA FA403 (.A(s_1_30_2), .B(s_2_30_2), .Cin(s_3_30_2), .S(s_2_30_1), .Cout(s_3_31_1));
    assign s_1_30_1 = s_4_30_2;
    FA FA404 (.A(s_1_31_2), .B(s_2_31_2), .Cin(s_3_31_2), .S(s_2_31_1), .Cout(s_3_32_1));
    assign s_1_31_1 = s_4_31_2;
    FA FA405 (.A(s_1_32_2), .B(s_2_32_2), .Cin(s_3_32_2), .S(s_2_32_1), .Cout(s_3_33_1));
    assign s_1_32_1 = s_4_32_2;
    // total 1 half adders and 28 full adders
    // d_2 = 3 done

    assign s_1_1_0 = s_1_1_1;
    assign s_2_2_0 = s_1_2_1;
    assign s_1_2_0 = s_2_2_1;
    HA HA29 (.A(s_1_3_1), .B(s_2_3_1), .S(s_2_3_0), .C(s_2_4_0));
    assign s_1_3_0 = s_3_3_1;
    FA FA406 (.A(s_1_4_1), .B(s_2_4_1), .Cin(s_3_4_1), .S(s_1_4_0), .Cout(s_2_5_0));
    FA FA407 (.A(s_1_5_1), .B(s_2_5_1), .Cin(s_3_5_1), .S(s_1_5_0), .Cout(s_2_6_0));
    FA FA408 (.A(s_1_6_1), .B(s_2_6_1), .Cin(s_3_6_1), .S(s_1_6_0), .Cout(s_2_7_0));
    FA FA409 (.A(s_1_7_1), .B(s_2_7_1), .Cin(s_3_7_1), .S(s_1_7_0), .Cout(s_2_8_0));
    FA FA410 (.A(s_1_8_1), .B(s_2_8_1), .Cin(s_3_8_1), .S(s_1_8_0), .Cout(s_2_9_0));
    FA FA411 (.A(s_1_9_1), .B(s_2_9_1), .Cin(s_3_9_1), .S(s_1_9_0), .Cout(s_2_10_0));
    FA FA412 (.A(s_1_10_1), .B(s_2_10_1), .Cin(s_3_10_1), .S(s_1_10_0), .Cout(s_2_11_0));
    FA FA413 (.A(s_1_11_1), .B(s_2_11_1), .Cin(s_3_11_1), .S(s_1_11_0), .Cout(s_2_12_0));
    FA FA414 (.A(s_1_12_1), .B(s_2_12_1), .Cin(s_3_12_1), .S(s_1_12_0), .Cout(s_2_13_0));
    FA FA415 (.A(s_1_13_1), .B(s_2_13_1), .Cin(s_3_13_1), .S(s_1_13_0), .Cout(s_2_14_0));
    FA FA416 (.A(s_1_14_1), .B(s_2_14_1), .Cin(s_3_14_1), .S(s_1_14_0), .Cout(s_2_15_0));
    FA FA417 (.A(s_1_15_1), .B(s_2_15_1), .Cin(s_3_15_1), .S(s_1_15_0), .Cout(s_2_16_0));
    FA FA418 (.A(s_1_16_1), .B(s_2_16_1), .Cin(s_3_16_1), .S(s_1_16_0), .Cout(s_2_17_0));
    FA FA419 (.A(s_1_17_1), .B(s_2_17_1), .Cin(s_3_17_1), .S(s_1_17_0), .Cout(s_2_18_0));
    FA FA420 (.A(s_1_18_1), .B(s_2_18_1), .Cin(s_3_18_1), .S(s_1_18_0), .Cout(s_2_19_0));
    FA FA421 (.A(s_1_19_1), .B(s_2_19_1), .Cin(s_3_19_1), .S(s_1_19_0), .Cout(s_2_20_0));
    FA FA422 (.A(s_1_20_1), .B(s_2_20_1), .Cin(s_3_20_1), .S(s_1_20_0), .Cout(s_2_21_0));
    FA FA423 (.A(s_1_21_1), .B(s_2_21_1), .Cin(s_3_21_1), .S(s_1_21_0), .Cout(s_2_22_0));
    FA FA424 (.A(s_1_22_1), .B(s_2_22_1), .Cin(s_3_22_1), .S(s_1_22_0), .Cout(s_2_23_0));
    FA FA425 (.A(s_1_23_1), .B(s_2_23_1), .Cin(s_3_23_1), .S(s_1_23_0), .Cout(s_2_24_0));
    FA FA426 (.A(s_1_24_1), .B(s_2_24_1), .Cin(s_3_24_1), .S(s_1_24_0), .Cout(s_2_25_0));
    FA FA427 (.A(s_1_25_1), .B(s_2_25_1), .Cin(s_3_25_1), .S(s_1_25_0), .Cout(s_2_26_0));
    FA FA428 (.A(s_1_26_1), .B(s_2_26_1), .Cin(s_3_26_1), .S(s_1_26_0), .Cout(s_2_27_0));
    FA FA429 (.A(s_1_27_1), .B(s_2_27_1), .Cin(s_3_27_1), .S(s_1_27_0), .Cout(s_2_28_0));
    FA FA430 (.A(s_1_28_1), .B(s_2_28_1), .Cin(s_3_28_1), .S(s_1_28_0), .Cout(s_2_29_0));
    FA FA431 (.A(s_1_29_1), .B(s_2_29_1), .Cin(s_3_29_1), .S(s_1_29_0), .Cout(s_2_30_0));
    FA FA432 (.A(s_1_30_1), .B(s_2_30_1), .Cin(s_3_30_1), .S(s_1_30_0), .Cout(s_2_31_0));
    FA FA433 (.A(s_1_31_1), .B(s_2_31_1), .Cin(s_3_31_1), .S(s_1_31_0), .Cout(s_2_32_0));
    FA FA434 (.A(s_1_32_1), .B(s_2_32_1), .Cin(s_3_32_1), .S(s_1_32_0), .Cout(s_2_33_0));
    // total 1 half adders and 29 full adders
    // d_1 = 2 done

    wire c_out_1, c_out_2, c_out_3, c_out_4, c_out_5, c_out_6, c_out_7, c_out_8, c_out_9, c_out_10, 
        c_out_11, c_out_12, c_out_13, c_out_14, c_out_15, c_out_16, c_out_17, c_out_18, c_out_19, c_out_20, 
        c_out_21, c_out_22, c_out_23, c_out_24, c_out_25, c_out_26, c_out_27, c_out_28, c_out_29, c_out_30, c_out_31;
    
    assign C[0] = s_1_1_0;
    HA HA30 (.A(s_1_2_0), .B(s_2_2_0), .S(C[1]), .C(c_out_1));
    FA FA435 (.A(s_1_3_0), .B(s_2_3_0), .Cin(c_out_1), .S(C[2]), .Cout(c_out_2));
    FA FA436 (.A(s_1_4_0), .B(s_2_4_0), .Cin(c_out_2), .S(C[3]), .Cout(c_out_3));
    FA FA437 (.A(s_1_5_0), .B(s_2_5_0), .Cin(c_out_3), .S(C[4]), .Cout(c_out_4));
    FA FA438 (.A(s_1_6_0), .B(s_2_6_0), .Cin(c_out_4), .S(C[5]), .Cout(c_out_5));
    FA FA439 (.A(s_1_7_0), .B(s_2_7_0), .Cin(c_out_5), .S(C[6]), .Cout(c_out_6));
    FA FA440 (.A(s_1_8_0), .B(s_2_8_0), .Cin(c_out_6), .S(C[7]), .Cout(c_out_7));
    FA FA441 (.A(s_1_9_0), .B(s_2_9_0), .Cin(c_out_7), .S(C[8]), .Cout(c_out_8));
    FA FA442 (.A(s_1_10_0), .B(s_2_10_0), .Cin(c_out_8), .S(C[9]), .Cout(c_out_9));
    FA FA443 (.A(s_1_11_0), .B(s_2_11_0), .Cin(c_out_9), .S(C[10]), .Cout(c_out_10));
    FA FA444 (.A(s_1_12_0), .B(s_2_12_0), .Cin(c_out_10), .S(C[11]), .Cout(c_out_11));
    FA FA445 (.A(s_1_13_0), .B(s_2_13_0), .Cin(c_out_11), .S(C[12]), .Cout(c_out_12));
    FA FA446 (.A(s_1_14_0), .B(s_2_14_0), .Cin(c_out_12), .S(C[13]), .Cout(c_out_13));
    FA FA447 (.A(s_1_15_0), .B(s_2_15_0), .Cin(c_out_13), .S(C[14]), .Cout(c_out_14));
    FA FA448 (.A(s_1_16_0), .B(s_2_16_0), .Cin(c_out_14), .S(C[15]), .Cout(c_out_15));
    FA FA449 (.A(s_1_17_0), .B(s_2_17_0), .Cin(c_out_15), .S(C[16]), .Cout(c_out_16));
    FA FA450 (.A(s_1_18_0), .B(s_2_18_0), .Cin(c_out_16), .S(C[17]), .Cout(c_out_17));
    FA FA451 (.A(s_1_19_0), .B(s_2_19_0), .Cin(c_out_17), .S(C[18]), .Cout(c_out_18));
    FA FA452 (.A(s_1_20_0), .B(s_2_20_0), .Cin(c_out_18), .S(C[19]), .Cout(c_out_19));
    FA FA453 (.A(s_1_21_0), .B(s_2_21_0), .Cin(c_out_19), .S(C[20]), .Cout(c_out_20));
    FA FA454 (.A(s_1_22_0), .B(s_2_22_0), .Cin(c_out_20), .S(C[21]), .Cout(c_out_21));
    FA FA455 (.A(s_1_23_0), .B(s_2_23_0), .Cin(c_out_21), .S(C[22]), .Cout(c_out_22));
    FA FA456 (.A(s_1_24_0), .B(s_2_24_0), .Cin(c_out_22), .S(C[23]), .Cout(c_out_23));
    FA FA457 (.A(s_1_25_0), .B(s_2_25_0), .Cin(c_out_23), .S(C[24]), .Cout(c_out_24));
    FA FA458 (.A(s_1_26_0), .B(s_2_26_0), .Cin(c_out_24), .S(C[25]), .Cout(c_out_25));
    FA FA459 (.A(s_1_27_0), .B(s_2_27_0), .Cin(c_out_25), .S(C[26]), .Cout(c_out_26));
    FA FA460 (.A(s_1_28_0), .B(s_2_28_0), .Cin(c_out_26), .S(C[27]), .Cout(c_out_27));
    FA FA461 (.A(s_1_29_0), .B(s_2_29_0), .Cin(c_out_27), .S(C[28]), .Cout(c_out_28));
    FA FA462 (.A(s_1_30_0), .B(s_2_30_0), .Cin(c_out_28), .S(C[29]), .Cout(c_out_29));
    FA FA463 (.A(s_1_31_0), .B(s_2_31_0), .Cin(c_out_29), .S(C[30]), .Cout(c_out_30));
    FA FA464 (.A(s_1_32_0), .B(s_2_32_0), .Cin(c_out_30), .S(C[31]), .Cout(c_out_31));

    // always@(posedge clk) begin
    //     if (~rst_n) begin
    //         A <= 0;
    //         B <= 0;
    //         C_r <= 0;
    //     end
    //     else begin
    //         A <= A;
    //         B <= B;
    //         C_r <= C;
    //     end
    // end

endmodule